-- fixed instruction memory
-- address : 15bit, capacity : 32Kwords
-- instruction length : 36bit
-- write only if opcode /= "100100"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity inst_mem_fixed is
  port (
    clk  : in  std_logic;
    addr : in  std_logic_vector(14 downto 0);
    din  : in  std_logic_vector(35 downto 0);
    inst : out std_logic_vector(35 downto 0);
    EN   : in  std_logic;
    WE   : in  std_logic);
end inst_mem_fixed;

architecture box of inst_mem_fixed is
  type mem_t is array(0 to 32767) of std_logic_vector(35 downto 0);
  signal mem : mem_t := (               -- 2nd_base/min_rt_2.s
"101001000000000111010000000110101100",--0
"101001000000000000010000000000000001",--1
"101000000001111000000001000000000000",--2
"001001000000000111010000000110101100",--3
"101001000000000111010000000110101010",--4
"001001111100000111110000000000000000",--5
"000111000000000000000111010110101010",--6
"101000000001111000000000100000000000",--7
"101110000001111000000001100000000000",--8
"101001000000000111010000000110101001",--9
"000111000000000000000111010110110001",--10
"001101000000000111010000000110101100",--11
"101000111011111000000001000000000000",--12
"101001111010000111010000000000001011",--13
"001001000100000000010000000000001010",--14
"001001000100000000010000000000001001",--15
"001001000100000000010000000000001000",--16
"001001000100000000010000000000000111",--17
"001001000100000000000000000000000110",--18
"001001000100000000010000000000000101",--19
"001001000100000000010000000000000100",--20
"001001000100000000000000000000000011",--21
"001001000100000000000000000000000010",--22
"001001000100000000000000000000000001",--23
"001001000100000000000000000000000000",--24
"001001000000000111010000000110101100",--25
"101001000000000111010000000101101101",--26
"101001000000000000010000000000111100",--27
"000111000000000000000111010110101010",--28
"101001000000000000010000000000000011",--29
"101110000001111000000001100000000000",--30
"101001000000000111010000000101101010",--31
"000111000000000000000111010110110001",--32
"101001000000000000010000000000000011",--33
"101110000001111000000001100000000000",--34
"101001000000000111010000000101100111",--35
"000111000000000000000111010110110001",--36
"101001000000000000010000000000000011",--37
"101110000001111000000001100000000000",--38
"101001000000000111010000000101100100",--39
"000111000000000000000111010110110001",--40
"101001000000000000010000000000000001",--41
"101111000001110000110100001101111111",--42
"101001000000000111010000000101100011",--43
"000111000000000000000111010110110001",--44
"001101111100000111110000000000000000",--45
"001101000000000111010000000110101100",--46
"101001000000000000010000000000110010",--47
"001001111100000000010000000000000000",--48
"101001000000000000010000000000000001",--49
"101001000000000000101111111111111111",--50
"001001111100000111111111111111111111",--51
"000111000000000000000111010110101010",--52
"101000000011111000000001000000000000",--53
"001001000000000111010000000110101100",--54
"101001000000000111010000000100110001",--55
"001101111100000000010000000000000000",--56
"000111000000000000000111010110101010",--57
"001101111100000111111111111111111111",--58
"001101000000000111010000000110101100",--59
"101001000000000000010000000000000001",--60
"001101000000000000100000000100110001",--61
"001001111100000000011111111111111111",--62
"101001000000000000010000000000000001",--63
"001001111100000111111111111111111110",--64
"000111000000000000000111010110101010",--65
"101000000011111000000001000000000000",--66
"001001000000000111010000000110101100",--67
"101001000000000111010000000100110000",--68
"001101111100000000011111111111111111",--69
"000111000000000000000111010110101010",--70
"101001000000000000010000000000000001",--71
"101110000001111000000001100000000000",--72
"101001000000000111010000000100101111",--73
"000111000000000000000111010110110001",--74
"101001000000000000010000000000000001",--75
"101000000001111000000001000000000000",--76
"101001000000000111010000000100101110",--77
"000111000000000000000111010110101010",--78
"101001000000000000010000000000000001",--79
"101111000111110000110100111001101110",--80
"101111000111100000110110101100101000",--81
"101001000000000111010000000100101101",--82
"000111000000000000000111010110110001",--83
"101001000000000000010000000000000011",--84
"101110000001111000000001100000000000",--85
"101001000000000111010000000100101010",--86
"000111000000000000000111010110110001",--87
"101001000000000000010000000000000001",--88
"101000000001111000000001000000000000",--89
"101001000000000111010000000100101001",--90
"000111000000000000000111010110101010",--91
"101001000000000000010000000000000011",--92
"101110000001111000000001100000000000",--93
"101001000000000111010000000100100110",--94
"000111000000000000000111010110110001",--95
"101001000000000000010000000000000011",--96
"101110000001111000000001100000000000",--97
"101001000000000111010000000100100011",--98
"000111000000000000000111010110110001",--99
"101001000000000000010000000000000011",--100
"101110000001111000000001100000000000",--101
"101001000000000111010000000100100000",--102
"000111000000000000000111010110110001",--103
"101001000000000000010000000000000011",--104
"101110000001111000000001100000000000",--105
"101001000000000111010000000100011101",--106
"000111000000000000000111010110110001",--107
"101001000000000000010000000000000010",--108
"101000000001111000000001000000000000",--109
"101001000000000111010000000100011011",--110
"000111000000000000000111010110101010",--111
"101001000000000000010000000000000010",--112
"101000000001111000000001000000000000",--113
"101001000000000111010000000100011001",--114
"000111000000000000000111010110101010",--115
"101001000000000000010000000000000001",--116
"101110000001111000000001100000000000",--117
"101001000000000111010000000100011000",--118
"000111000000000000000111010110110001",--119
"101001000000000000010000000000000011",--120
"101110000001111000000001100000000000",--121
"101001000000000111010000000100010101",--122
"000111000000000000000111010110110001",--123
"101001000000000000010000000000000011",--124
"101110000001111000000001100000000000",--125
"101001000000000111010000000100010010",--126
"000111000000000000000111010110110001",--127
"101001000000000000010000000000000011",--128
"101110000001111000000001100000000000",--129
"101001000000000111010000000100001111",--130
"000111000000000000000111010110110001",--131
"101001000000000000010000000000000011",--132
"101110000001111000000001100000000000",--133
"101001000000000111010000000100001100",--134
"000111000000000000000111010110110001",--135
"101001000000000000010000000000000011",--136
"101110000001111000000001100000000000",--137
"101001000000000111010000000100001001",--138
"000111000000000000000111010110110001",--139
"101001000000000000010000000000000011",--140
"101110000001111000000001100000000000",--141
"101001000000000111010000000100000110",--142
"000111000000000000000111010110110001",--143
"101000000001111000000000100000000000",--144
"101110000001111000000001100000000000",--145
"101001000000000111010000000100000101",--146
"000111000000000000000111010110110001",--147
"001101111100000111111111111111111110",--148
"101001000000000111010000000100000100",--149
"001001111100000000011111111111111110",--150
"101000000001111000000000100000000000",--151
"101001000000000000100000000100000101",--152
"001001111100000111111111111111111101",--153
"000111000000000000000111010110101010",--154
"001101000000000111010000000110101100",--155
"101000111011111000000001000000000000",--156
"101001111010000111010000000000000010",--157
"001001000100000000010000000000000001",--158
"001101111100000000011111111111111110",--159
"001001000100000000010000000000000000",--160
"001001000000000111010000000110101100",--161
"101001000000000111010000000100000011",--162
"101000000001111000000000100000000000",--163
"000111000000000000000111010110101010",--164
"101001000000000000010000000000000101",--165
"101001000000000111010000000011111110",--166
"101001000000000000100000000100000011",--167
"000111000000000000000111010110101010",--168
"101000000001111000000000100000000000",--169
"101110000001111000000001100000000000",--170
"101001000000000111010000000011111101",--171
"000111000000000000000111010110110001",--172
"101001000000000000010000000000000011",--173
"101110000001111000000001100000000000",--174
"101001000000000111010000000011111010",--175
"000111000000000000000111010110110001",--176
"001101111100000111111111111111111101",--177
"101001000000000111010000000010111110",--178
"001001111100000000011111111111111101",--179
"101001000000000000010000000000111100",--180
"101001000000000000100000000011111101",--181
"001001111100000111111111111111111100",--182
"000111000000000000000111010110101010",--183
"001001000000000000010000000010111101",--184
"001101111100000000011111111111111101",--185
"001001000000000000010000000010111100",--186
"101000000001111000000000100000000000",--187
"101110000001111000000001100000000000",--188
"101001000000000111010000000010111011",--189
"000111000000000000000111010110110001",--190
"001101111100000111111111111111111100",--191
"101001000000000111010000000010111010",--192
"001001111100000000011111111111111100",--193
"101000000001111000000000100000000000",--194
"101001000000000000100000000010111011",--195
"001001111100000111111111111111111011",--196
"000111000000000000000111010110101010",--197
"001001000000000000010000000010111001",--198
"001101111100000000011111111111111100",--199
"001001000000000000010000000010111000",--200
"101001000000000000010000000010111000",--201
"001101000000000111010000000110101100",--202
"101000111011111000000001000000000000",--203
"101001111010000111010000000000000011",--204
"001011000100000000000000000000000010",--205
"001001000100000000010000000000000001",--206
"001001000100000000000000000000000000",--207
"001001000000000111010000000110101100",--208
"101001000000000111010000000000000100",--209
"101001000000000000010000000010110100",--210
"000111000000000000000111010110101010",--211
"101001000000000000010000000000000001",--212
"101000000001111000000001000000000000",--213
"101001000000000111010000000000000011",--214
"000111000000000000000111010110101010",--215
"001101000000000111010000000110101100",--216
"101001000000000000010000000000000010",--217
"101001000000000000100000000000000010",--218
"001001000000000000010000000100011011",--219
"001001000000000000100000000100011100",--220
"101001000000000000100000000000000001",--221
"001001000000000000100000000100011001",--222
"101001000000000000100000000000000001",--223
"001001000000000000100000000100011010",--224
"101111000001110000110100001100000000",--225
"101010000011101000000010000000000000",--226
"111110001000011000000010000000000000",--227
"111110000110001001000001100000000000",--228
"001011000000000000110000000100011000",--229
"101001111100010111100000000000000110",--230
"000111000000000000000110101111000000",--231
"101001111100000111100000000000000110",--232
"001101111100000111111111111111111011",--233
"001001000000000000010000000000000010",--234
"001001111100000000011111111111111011",--235
"001001111100000111111111111111111010",--236
"101001111100010111100000000000000111",--237
"000111000000000000000110101111000000",--238
"101001111100000111100000000000000111",--239
"001101111100000111111111111111111010",--240
"001001000000000000010000000000000001",--241
"001001111100000000011111111111111010",--242
"001001111100000111111111111111111001",--243
"101001111100010111100000000000001000",--244
"000111000000000000000110101111000000",--245
"101001111100000111100000000000001000",--246
"001101111100000111111111111111111001",--247
"001001000000000000010000000000000000",--248
"000011000000000000000001100000000000",--249
"001011000000000000110000000101101010",--250
"000011000000000000000001100000000000",--251
"001011000000000000110000000101101011",--252
"000011000000000000000001100000000000",--253
"001011000000000000110000000101101100",--254
"000011000000000000000001100000000000",--255
"101111001001110001000011110010001110",--256
"101111001001100001001111101000110101",--257
"111110000110001001000001100000000000",--258
"001001111100000000011111111111111001",--259
"001011111100000000111111111111111000",--260
"001001111100000111111111111111110111",--261
"000111000000000000000111010110111000",--262
"001101111100000111111111111111110111",--263
"001111111100000001001111111111111000",--264
"001011111100000000111111111111110111",--265
"101110001001111000000001100000000000",--266
"001001111100000111111111111111110110",--267
"000111000000000000000111011000000010",--268
"001101111100000111111111111111110110",--269
"000011000000000000000010000000000000",--270
"101111001011110001010011110010001110",--271
"101111001011100001011111101000110101",--272
"111110001000001001010010000000000000",--273
"001011111100000000111111111111110110",--274
"001011111100000001001111111111110101",--275
"101110001001111000000001100000000000",--276
"001001111100000111111111111111110100",--277
"000111000000000000000111010110111000",--278
"001101111100000111111111111111110100",--279
"001111111100000001001111111111110101",--280
"001011111100000000111111111111110100",--281
"101110001001111000000001100000000000",--282
"001001111100000111111111111111110011",--283
"000111000000000000000111011000000010",--284
"001101111100000111111111111111110011",--285
"001111111100000001001111111111110111",--286
"111110001000001000110010100000000000",--287
"101111000001110001100100001101001000",--288
"111110001010001001100010100000000000",--289
"001011000000000001010000000100001001",--290
"101111000001110001011100001101001000",--291
"001111111100000001101111111111110110",--292
"111110001100001001010010100000000000",--293
"001011000000000001010000000100001010",--294
"001111111100000001011111111111110100",--295
"111110001000001001010011100000000000",--296
"101111000001110010000100001101001000",--297
"111110001110001010000011100000000000",--298
"001011000000000001110000000100001011",--299
"001011000000000001010000000100001111",--300
"001011000000000000000000000100010000",--301
"101110000111111000000011100000000010",--302
"001011000000000001110000000100010001",--303
"101110001101111000000011100000000010",--304
"111110001110001000110001100000000000",--305
"001011000000000000110000000100001100",--306
"101110001001111000000001100000000010",--307
"001011000000000000110000000100001101",--308
"111110001100001001010001100000000010",--309
"001011000000000000110000000100001110",--310
"001111000000000000110000000101101010",--311
"001111000000000001000000000100001001",--312
"111110000110010001000001100000000000",--313
"001011000000000000110000000101100111",--314
"001111000000000000110000000101101011",--315
"001111000000000001000000000100001010",--316
"111110000110010001000001100000000000",--317
"001011000000000000110000000101101000",--318
"001111000000000000110000000101101100",--319
"001111000000000001000000000100001011",--320
"111110000110010001000001100000000000",--321
"001011000000000000110000000101101001",--322
"000010000000000000000000100000000000",--323
"000011000000000000000001100000000000",--324
"101111001001110001000011110010001110",--325
"101111001001100001001111101000110101",--326
"111110000110001001000001100000000000",--327
"001011111100000000111111111111110011",--328
"001001111100000111111111111111110010",--329
"000111000000000000000111011000000010",--330
"001101111100000111111111111111110010",--331
"101110000111111000000001100000000010",--332
"001011000000000000110000000101100101",--333
"000011000000000000000001100000000000",--334
"101111001001110001000011110010001110",--335
"101111001001100001001111101000110101",--336
"111110000110001001000001100000000000",--337
"001111111100000001001111111111110011",--338
"001011111100000000111111111111110010",--339
"101110001001111000000001100000000000",--340
"001001111100000111111111111111110001",--341
"000111000000000000000111010110111000",--342
"001101111100000111111111111111110001",--343
"001111111100000001001111111111110010",--344
"001011111100000000111111111111110001",--345
"101110001001111000000001100000000000",--346
"001001111100000111111111111111110000",--347
"000111000000000000000111011000000010",--348
"001111111100000001001111111111110001",--349
"111110001000001000110001100000000000",--350
"001011000000000000110000000101100100",--351
"001111111100000000111111111111110010",--352
"000111000000000000000111010110111000",--353
"001111111100000001001111111111110001",--354
"111110001000001000110001100000000000",--355
"001011000000000000110000000101100110",--356
"000011000000000000000001100000000000",--357
"001011000000000000110000000101100011",--358
"101000000001111000000000100000000000",--359
"101001111100010111100000000000010001",--360
"000111000000000000000000010000000001",--361
"101001111100000111100000000000010001",--362
"101000000001111000000000100000000000",--363
"101001111100010111100000000000010001",--364
"000111000000000000000000010101111100",--365
"101001111100000111100000000000010001",--366
"101000000001111000000000100000000000",--367
"101001111100010111100000000000010001",--368
"000111000000000000000000010101100011",--369
"101001111100000111100000000000010001",--370
"001101111100000111111111111111110000",--371
"001001000000000000010000000100110000",--372
"101001000000000000010000000001010000",--373
"000000000010000000000000000000000000",--374
"101001000000000000010000000000110110",--375
"000000000010000000000000000000000000",--376
"101001000000000000010000000000001010",--377
"000000000010000000000000000000000000",--378
"001101000000000000010000000100011011",--379
"011011000011011001000000000000000010",--380
"101000000001111000000001000000000000",--381
"000101000000000000000000000110011111",--382
"011011000011110010000000000000000010",--383
"101001000000000000100000000000000001",--384
"000101000000000000000000000110011111",--385
"101001000000000000100000000100101100",--386
"010100000101000000010000000000000010",--387
"101001000000000000100000000000000010",--388
"000101000000000000000000000110011111",--389
"101001000000000000100000000110010000",--390
"010100000101000000010000000000000010",--391
"101001000000000000100000000000000011",--392
"000101000000000000000000000110011111",--393
"101001000000000000100000000111110100",--394
"010100000101000000010000000000000010",--395
"101001000000000000100000000000000100",--396
"000101000000000000000000000110011111",--397
"101001000000000000100000001001011000",--398
"010100000101000000010000000000000010",--399
"101001000000000000100000000000000101",--400
"000101000000000000000000000110011111",--401
"101001000000000000100000001010111100",--402
"010100000101000000010000000000000010",--403
"101001000000000000100000000000000110",--404
"000101000000000000000000000110011111",--405
"101001000000000000100000001100100000",--406
"010100000101000000010000000000000010",--407
"101001000000000000100000000000000111",--408
"000101000000000000000000000110011111",--409
"101001000000000000100000001110000100",--410
"010100000101000000010000000000000010",--411
"101001000000000000100000000000001000",--412
"000101000000000000000000000110011111",--413
"101001000000000000100000000000001001",--414
"101000000101000000110001100110000110",--415
"101000000101000001000010000101000101",--416
"101000000110000001000001100000000000",--417
"101000000101000001000010000010000010",--418
"101000000110000001000001100000000000",--419
"101000000010010000110000100000000000",--420
"011011000011000010100000000000000010",--421
"101000000001111000000001100000000000",--422
"000101000000000000000000000111000001",--423
"011011000011000101000000000000000010",--424
"101001000000000000110000000000000001",--425
"000101000000000000000000000111000001",--426
"011011000011000111100000000000000010",--427
"101001000000000000110000000000000010",--428
"000101000000000000000000000111000001",--429
"011011000011001010000000000000000010",--430
"101001000000000000110000000000000011",--431
"000101000000000000000000000111000001",--432
"011011000011001100100000000000000010",--433
"101001000000000000110000000000000100",--434
"000101000000000000000000000111000001",--435
"011011000011001111000000000000000010",--436
"101001000000000000110000000000000101",--437
"000101000000000000000000000111000001",--438
"011011000011010001100000000000000010",--439
"101001000000000000110000000000000110",--440
"000101000000000000000000000111000001",--441
"011011000011010100000000000000000010",--442
"101001000000000000110000000000000111",--443
"000101000000000000000000000111000001",--444
"011011000011010110100000000000000010",--445
"101001000000000000110000000000001000",--446
"000101000000000000000000000111000001",--447
"101001000000000000110000000000001001",--448
"101000000111000001000010000011000011",--449
"101000000111000001010010100001000001",--450
"101000001000000001010010000000000000",--451
"101000000010010001000000100000000000",--452
"011100000101000000000000000000001001",--453
"011100000111000000000000000000000011",--454
"101001000010000000010000000000110000",--455
"000000000010000000000000000000000000",--456
"000101000000000000000000000111010101",--457
"101001000110000000100000000000110000",--458
"000000000100000000000000000000000000",--459
"101001000010000000010000000000110000",--460
"000000000010000000000000000000000000",--461
"000101000000000000000000000111010101",--462
"101001000100000000100000000000110000",--463
"000000000100000000000000000000000000",--464
"101001000110000000100000000000110000",--465
"000000000100000000000000000000000000",--466
"101001000010000000010000000000110000",--467
"000000000010000000000000000000000000",--468
"101001000000000000010000000000100000",--469
"000000000010000000000000000000000000",--470
"001101000000000000010000000100011100",--471
"011011000011011001000000000000000010",--472
"101000000001111000000001000000000000",--473
"000101000000000000000000000111111011",--474
"011011000011110010000000000000000010",--475
"101001000000000000100000000000000001",--476
"000101000000000000000000000111111011",--477
"101001000000000000100000000100101100",--478
"010100000101000000010000000000000010",--479
"101001000000000000100000000000000010",--480
"000101000000000000000000000111111011",--481
"101001000000000000100000000110010000",--482
"010100000101000000010000000000000010",--483
"101001000000000000100000000000000011",--484
"000101000000000000000000000111111011",--485
"101001000000000000100000000111110100",--486
"010100000101000000010000000000000010",--487
"101001000000000000100000000000000100",--488
"000101000000000000000000000111111011",--489
"101001000000000000100000001001011000",--490
"010100000101000000010000000000000010",--491
"101001000000000000100000000000000101",--492
"000101000000000000000000000111111011",--493
"101001000000000000100000001010111100",--494
"010100000101000000010000000000000010",--495
"101001000000000000100000000000000110",--496
"000101000000000000000000000111111011",--497
"101001000000000000100000001100100000",--498
"010100000101000000010000000000000010",--499
"101001000000000000100000000000000111",--500
"000101000000000000000000000111111011",--501
"101001000000000000100000001110000100",--502
"010100000101000000010000000000000010",--503
"101001000000000000100000000000001000",--504
"000101000000000000000000000111111011",--505
"101001000000000000100000000000001001",--506
"101000000101000000110001100110000110",--507
"101000000101000001000010000101000101",--508
"101000000110000001000001100000000000",--509
"101000000101000001000010000010000010",--510
"101000000110000001000001100000000000",--511
"101000000010010000110000100000000000",--512
"011011000011000010100000000000000010",--513
"101000000001111000000001100000000000",--514
"000101000000000000000000001000011101",--515
"011011000011000101000000000000000010",--516
"101001000000000000110000000000000001",--517
"000101000000000000000000001000011101",--518
"011011000011000111100000000000000010",--519
"101001000000000000110000000000000010",--520
"000101000000000000000000001000011101",--521
"011011000011001010000000000000000010",--522
"101001000000000000110000000000000011",--523
"000101000000000000000000001000011101",--524
"011011000011001100100000000000000010",--525
"101001000000000000110000000000000100",--526
"000101000000000000000000001000011101",--527
"011011000011001111000000000000000010",--528
"101001000000000000110000000000000101",--529
"000101000000000000000000001000011101",--530
"011011000011010001100000000000000010",--531
"101001000000000000110000000000000110",--532
"000101000000000000000000001000011101",--533
"011011000011010100000000000000000010",--534
"101001000000000000110000000000000111",--535
"000101000000000000000000001000011101",--536
"011011000011010110100000000000000010",--537
"101001000000000000110000000000001000",--538
"000101000000000000000000001000011101",--539
"101001000000000000110000000000001001",--540
"101000000111000001000010000011000011",--541
"101000000111000001010010100001000001",--542
"101000001000000001010010000000000000",--543
"101000000010010001000000100000000000",--544
"011100000101000000000000000000001001",--545
"011100000111000000000000000000000011",--546
"101001000010000000010000000000110000",--547
"000000000010000000000000000000000000",--548
"000101000000000000000000001000110001",--549
"101001000110000000100000000000110000",--550
"000000000100000000000000000000000000",--551
"101001000010000000010000000000110000",--552
"000000000010000000000000000000000000",--553
"000101000000000000000000001000110001",--554
"101001000100000000100000000000110000",--555
"000000000100000000000000000000000000",--556
"101001000110000000100000000000110000",--557
"000000000100000000000000000000000000",--558
"101001000010000000010000000000110000",--559
"000000000010000000000000000000000000",--560
"101001000000000000010000000000100000",--561
"000000000010000000000000000000000000",--562
"101001000000000000010000000000110010",--563
"000000000010000000000000000000000000",--564
"101001000000000000010000000000110101",--565
"000000000010000000000000000000000000",--566
"101001000000000000010000000000110101",--567
"000000000010000000000000000000000000",--568
"101001000000000000010000000000001010",--569
"000000000010000000000000000000000000",--570
"101001000000000000010000000000000100",--571
"001001111100000111111111111111110000",--572
"101001111100010111100000000000010001",--573
"000111000000000000000111010100111111",--574
"101001111100000111100000000000010001",--575
"101001000000000000010000000000001001",--576
"101000000001111000000001000000000000",--577
"101000000001111000000001100000000000",--578
"101010000011101000000001100000000000",--579
"101111001001110001000011111001001100",--580
"101111001001100001001100110011001101",--581
"111110000110001001000001100000000000",--582
"101111001001110001000011111101100110",--583
"101111001001100001000110011001100110",--584
"111110000110010001000001100000000000",--585
"101001000000000000010000000000000100",--586
"101001111100010111100000000000010001",--587
"000111000000000000000110111011001001",--588
"101001111100000111100000000000010001",--589
"101001000000000000010000000000001000",--590
"101001000000000000100000000000000010",--591
"101001000000000000110000000000000100",--592
"101001111100010111100000000000010001",--593
"000111000000000000000111001001010001",--594
"101001111100000111100000000000010001",--595
"101001000000000000010000000000000100",--596
"101001111100010111100000000000010001",--597
"000111000000000000000111010101101110",--598
"101001111100000111100000000000010001",--599
"001111000000000000110000000101100100",--600
"001011000000000000110000000011111010",--601
"001111000000000000110000000101100101",--602
"001011000000000000110000000011111011",--603
"001111000000000000110000000101100110",--604
"001011000000000000110000000011111100",--605
"101001000000000000010000000010111100",--606
"101001111100010111100000000000010001",--607
"000111000000000000000000011001101010",--608
"101001111100000111100000000000010001",--609
"001101111100000111111111111111110000",--610
"001101000000000000010000000110101010",--611
"101001000010010000010000000000000001",--612
"010111000011000000000000000001101011",--613
"001101000010000000100000000101101101",--614
"001101000100000000110000000000000010",--615
"011111000111000000100000000001101000",--616
"001101000100000000110000000000000111",--617
"001111000110000000110000000000000000",--618
"011010000111000000010000000001100101",--619
"001101000100000001000000000000000001",--620
"011111001001000000010000000000110000",--621
"101000000011000000010000100010000010",--622
"001101000000000000100000000000000011",--623
"111110000110010000010001100000000010",--624
"001111000000010001000000000101100100",--625
"001111000000010001010000000101100101",--626
"001111000000010001100000000101100110",--627
"101001000010000000110000000000000001",--628
"001111000000000001110000000101100100",--629
"001011111100000001011111111111110000",--630
"001011111100000001101111111111101111",--631
"001011111100000001001111111111101110",--632
"001011111100000000111111111111101101",--633
"001001111100000000011111111111101100",--634
"001001111100000000101111111111101011",--635
"101000000101111000000000100000000000",--636
"101000000111111000000001000000000000",--637
"101110001111111000000010000000000000",--638
"001001111100000111111111111111101010",--639
"101001111100010111100000000000010111",--640
"000111000000000000000111010101111100",--641
"101001111100000111100000000000010111",--642
"001101111100000000011111111111101011",--643
"101001000010000000010000000000000001",--644
"001101111100000000111111111111101100",--645
"101001000110000000100000000000000010",--646
"001111000000000001010000000101100101",--647
"001111111100000000111111111111101101",--648
"001111111100000001001111111111101110",--649
"001111111100000001101111111111101111",--650
"101001111100010111100000000000010111",--651
"000111000000000000000111010101111100",--652
"101001111100000111100000000000010111",--653
"001101111100000000011111111111101011",--654
"101001000010000000010000000000000010",--655
"001101111100000000111111111111101100",--656
"101001000110000000100000000000000011",--657
"001111000000000001100000000101100110",--658
"001111111100000000111111111111101101",--659
"001111111100000001001111111111101110",--660
"001111111100000001011111111111110000",--661
"101001111100010111100000000000010111",--662
"000111000000000000000111010101111100",--663
"101001111100000111100000000000010111",--664
"001101111100000111111111111111101010",--665
"001101111100000000011111111111101011",--666
"101001000010000000010000000000000011",--667
"001001000000000000010000000000000011",--668
"000101000000000000000000001011010001",--669
"011111001001000000100000000000110010",--670
"101000000011000000010000100010000010",--671
"101001000010000000010000000000000001",--672
"001101000000000001000000000000000011",--673
"001111000110000000110000000000000000",--674
"111110000110010000010001100000000010",--675
"001101000100000000100000000000000100",--676
"001111000000000001000000000101100100",--677
"001111000100000001010000000000000000",--678
"111110001000001001010010000000000000",--679
"001111000000000001010000000101100101",--680
"001111000100000001100000000000000001",--681
"111110001010001001100010100000000000",--682
"111110001000000001010010000000000000",--683
"001111000000000001010000000101100110",--684
"001111000100000001100000000000000010",--685
"111110001010001001100010100000000000",--686
"111110001000000001010010000000000000",--687
"101111000001110001010100000000000000",--688
"001111000100000001100000000000000000",--689
"111110001010001001100010100000000000",--690
"111110001010001001000010100000000000",--691
"001111000000000001100000000101100100",--692
"111110001010010001100010100000000000",--693
"101111000001110001100100000000000000",--694
"001111000100000001110000000000000001",--695
"111110001100001001110011000000000000",--696
"111110001100001001000011000000000000",--697
"001111000000000001110000000101100101",--698
"111110001100010001110011000000000000",--699
"101111000001110001110100000000000000",--700
"001111000100000010000000000000000010",--701
"111110001110001010000011100000000000",--702
"111110001110001001000010000000000000",--703
"001111000000000001110000000101100110",--704
"111110001000010001110010000000000000",--705
"001001111100000001001111111111110000",--706
"101000000011111000000001000000000000",--707
"101000001001111000000000100000000000",--708
"101110001101111000001111100000000000",--709
"101110001001111000000011000000000000",--710
"101110001011111000000010000000000000",--711
"101110111111111000000010100000000000",--712
"001001111100000111111111111111101111",--713
"101001111100010111100000000000010010",--714
"000111000000000000000111010101111100",--715
"101001111100000111100000000000010010",--716
"001101111100000111111111111111101111",--717
"001101111100000000011111111111110000",--718
"101001000010000000010000000000000001",--719
"001001000000000000010000000000000011",--720
"001101000000000000010000000100011011",--721
"101001000010010000010000000000000001",--722
"010111000011000000000000000001101111",--723
"101000000001111000000001000000000000",--724
"001111000000000000110000000100011000",--725
"001101000000000000110000000100011010",--726
"101000000000010000110001100000000000",--727
"101010000111101000000010000000000000",--728
"111110000110001001000001100000000000",--729
"001111000000000001000000000100001100",--730
"111110000110001001000010000000000000",--731
"001111000000000001010000000100001001",--732
"111110001000000001010010000000000000",--733
"001111000000000001010000000100001101",--734
"111110000110001001010010100000000000",--735
"001111000000000001100000000100001010",--736
"111110001010000001100010100000000000",--737
"001111000000000001100000000100001110",--738
"111110000110001001100001100000000000",--739
"001111000000000001100000000100001011",--740
"111110000110000001100001100000000000",--741
"001111000000000001100000000100011000",--742
"001101000000000000110000000100011001",--743
"101000000010010000110001100000000000",--744
"101010000111101000000011100000000000",--745
"111110001100001001110011000000000000",--746
"001111000000000001110000000100001111",--747
"111110001100001001110011100000000000",--748
"111110001110000001000011100000000000",--749
"001011000000000001110000000100000110",--750
"001111000000000001110000000100010000",--751
"111110001100001001110011100000000000",--752
"111110001110000001010011100000000000",--753
"001011000000000001110000000100000111",--754
"001111000000000001110000000100010001",--755
"111110001100001001110011000000000000",--756
"111110001100000000110011000000000000",--757
"001011000000000001100000000100001000",--758
"001111000000000001100000000100000110",--759
"111110001100001001100011000000000000",--760
"001111000000000001110000000100000111",--761
"111110001110001001110011100000000000",--762
"111110001100000001110011000000000000",--763
"001111000000000001110000000100001000",--764
"111110001110001001110011100000000000",--765
"111110001100000001110011000000000000",--766
"111110001100100000000011000000000000",--767
"011110001101000000000000000000000010",--768
"101110000011111000000011000000000000",--769
"000101000000000000000000001100000100",--770
"111110001100011000000011000000000000",--771
"001111000000000001110000000100000110",--772
"111110001110001001100011100000000000",--773
"001011000000000001110000000100000110",--774
"001111000000000001110000000100000111",--775
"111110001110001001100011100000000000",--776
"001011000000000001110000000100000111",--777
"001111000000000001110000000100001000",--778
"111110001110001001100011000000000000",--779
"001011000000000001100000000100001000",--780
"001011000000000000000000000100011101",--781
"001011000000000000000000000100011110",--782
"001011000000000000000000000100011111",--783
"001111000000000001100000000101100111",--784
"001011000000000001100000000100010101",--785
"001111000000000001100000000101101000",--786
"001011000000000001100000000100010110",--787
"001111000000000001100000000101101001",--788
"001011000000000001100000000100010111",--789
"001101111100000001011111111111111010",--790
"001100001010000000010001100000000000",--791
"001011111100000000111111111111110000",--792
"001011111100000001011111111111101111",--793
"001011111100000001001111111111101110",--794
"001001111100000000101111111111101101",--795
"001001111100000000011111111111101100",--796
"101001000000000000100000000100000110",--797
"101000000001111000000000100000000000",--798
"101110000001111000000010000000000000",--799
"101110000011111000000001100000000000",--800
"001001111100000111111111111111101011",--801
"101001111100010111100000000000010110",--802
"000111000000000000000011010111001111",--803
"101001111100000111100000000000010110",--804
"001101111100000000011111111111101100",--805
"001101111100000000111111111111111010",--806
"001100000110000000010001000000000000",--807
"001101000100000000100000000000000000",--808
"001111000000000000110000000100011101",--809
"001011000100000000110000000000000000",--810
"001111000000000000110000000100011110",--811
"001011000100000000110000000000000001",--812
"001111000000000000110000000100011111",--813
"001011000100000000110000000000000010",--814
"001100000110000000010001000000000000",--815
"001101000100000000100000000000000110",--816
"001101111100000001001111111111101101",--817
"001001000100000001000000000000000000",--818
"001100000110000000010000100000000000",--819
"101000000001111000000001000000000000",--820
"101001111100010111100000000000010110",--821
"000111000000000000000110001000010000",--822
"101001111100000111100000000000010110",--823
"001101111100000000011111111111101100",--824
"101001000010010000100000000000000001",--825
"101001000000000000110000000000000001",--826
"001111111100000000111111111111101110",--827
"001111111100000001001111111111101111",--828
"001111111100000001011111111111110000",--829
"001101111100000000011111111111111010",--830
"101001111100010111100000000000010110",--831
"000111000000000000000110010100111001",--832
"101001111100000111100000000000010110",--833
"001101111100000111111111111111101011",--834
"101000000001111000000000100000000000",--835
"101001000000000001010000000000000010",--836
"001101111100000000101111111111111011",--837
"001101111100000000111111111111111010",--838
"001101111100000001001111111111111001",--839
"001001111100000111111111111111110000",--840
"101001111100010111100000000000010001",--841
"000111000000000000000110101011011010",--842
"100111000000000000000000000000000000",--843
"101111000001110001100011111100000000",--844
"010110001101000000110000000000000010",--845
"101110001011111000000001100000000000",--846
"000100000000000000001111100000000000",--847
"111110000110010000010011000000000000",--848
"111110000110001000110011100000000000",--849
"111110001110001001000011100000000000",--850
"111110000110000000110001100000000000",--851
"111110000110000000010001100000000000",--852
"111110000110000001010001100000000000",--853
"111110000110011000000001100000000000",--854
"111110001110001000110001100000000000",--855
"101111000001110001010011111100000000",--856
"010110001011000001100000000000000001",--857
"000100000000000000001111100000000000",--858
"111110001100010000010010100000000000",--859
"111110001100001001100011100000000000",--860
"111110001110001001000011100000000000",--861
"111110001100000001100011000000000000",--862
"111110001100000000010011000000000000",--863
"111110001100000000110001100000000000",--864
"111110000110011000000001100000000000",--865
"111110001110001000110001100000000000",--866
"101111000001110001100011111100000000",--867
"010110001101000001010000000000000001",--868
"000100000000000000001111100000000000",--869
"111110001010010000010011000000000000",--870
"111110001010001001010011100000000000",--871
"111110001110001001000011100000000000",--872
"111110001010000001010010100000000000",--873
"111110001010000000010010100000000000",--874
"111110001010000000110001100000000000",--875
"111110000110011000000001100000000000",--876
"111110001110001000110001100000000000",--877
"101111000001110001010011111100000000",--878
"010110001011000001100000000000000001",--879
"000100000000000000001111100000000000",--880
"111110001100010000010010100000000000",--881
"111110001100001001100011100000000000",--882
"111110001110001001000011100000000000",--883
"111110001100000001100011000000000000",--884
"111110001100000000010011000000000000",--885
"111110001100000000110001100000000000",--886
"111110000110011000000001100000000000",--887
"111110001110001000110001100000000000",--888
"101111000001110001100011111100000000",--889
"010110001101000001010000000000000001",--890
"000100000000000000001111100000000000",--891
"111110001010010000010011000000000000",--892
"111110001010001001010011100000000000",--893
"111110001110001001000011100000000000",--894
"111110001010000001010010100000000000",--895
"111110001010000000010010100000000000",--896
"111110001010000000110001100000000000",--897
"111110000110011000000001100000000000",--898
"111110001110001000110001100000000000",--899
"101111000001110001010011111100000000",--900
"010110001011000001100000000000000001",--901
"000100000000000000001111100000000000",--902
"111110001100010000010010100000000000",--903
"111110001100001001100011100000000000",--904
"111110001110001001000011100000000000",--905
"111110001100000001100011000000000000",--906
"111110001100000000010011000000000000",--907
"111110001100000000110001100000000000",--908
"111110000110011000000001100000000000",--909
"111110001110001000110001100000000000",--910
"101111000001110001100011111100000000",--911
"010110001101000001010000000000000001",--912
"000100000000000000001111100000000000",--913
"111110001010010000010011000000000000",--914
"111110001010001001010011100000000000",--915
"111110001110001001000011100000000000",--916
"111110001010000001010010100000000000",--917
"111110001010000000010010100000000000",--918
"111110001010000000110001100000000000",--919
"111110000110011000000001100000000000",--920
"111110001110001000110001100000000000",--921
"101111000001110001010011111100000000",--922
"010110001011000001100000000000000001",--923
"000100000000000000001111100000000000",--924
"111110001100010000010010100000000000",--925
"111110001100001001100011100000000000",--926
"111110001110001001000011100000000000",--927
"111110001100000001100011000000000000",--928
"111110001100000000010011000000000000",--929
"111110001100000000110001100000000000",--930
"111110000110011000000001100000000000",--931
"111110001110001000110001100000000000",--932
"101111000001110001100011111100000000",--933
"010110001101000001010000000000000001",--934
"000100000000000000001111100000000000",--935
"111110001010010000010011000000000000",--936
"111110001010001001010011100000000000",--937
"111110001110001001000011100000000000",--938
"111110001010000001010010100000000000",--939
"111110001010000000010010100000000000",--940
"111110001010000000110001100000000000",--941
"111110000110011000000001100000000000",--942
"111110001110001000110001100000000000",--943
"101111000001110001010011111100000000",--944
"010110001011000001100000000000000001",--945
"000100000000000000001111100000000000",--946
"111110001100010000010010100000000000",--947
"111110001100001001100011100000000000",--948
"111110001110001001000011100000000000",--949
"111110001100000001100011000000000000",--950
"111110001100000000010011000000000000",--951
"111110001100000000110001100000000000",--952
"111110000110011000000001100000000000",--953
"111110001110001000110001100000000000",--954
"101111000001110001100011111100000000",--955
"010110001101000001010000000000000001",--956
"000100000000000000001111100000000000",--957
"111110001010010000010011000000000000",--958
"111110001010001001010011100000000000",--959
"111110001110001001000011100000000000",--960
"111110001010000001010010100000000000",--961
"111110001010000000010010100000000000",--962
"111110001010000000110001100000000000",--963
"111110000110011000000001100000000000",--964
"111110001110001000110001100000000000",--965
"101111000001110001010011111100000000",--966
"010110001011000001100000000000000001",--967
"000100000000000000001111100000000000",--968
"111110001100010000010010100000000000",--969
"111110001100001001100011100000000000",--970
"111110001110001001000011100000000000",--971
"111110001100000001100011000000000000",--972
"111110001100000000010011000000000000",--973
"111110001100000000110001100000000000",--974
"111110000110011000000001100000000000",--975
"111110001110001000110001100000000000",--976
"101111000001110001100011111100000000",--977
"010110001101000001010000000000000001",--978
"000100000000000000001111100000000000",--979
"111110001010010000010011000000000000",--980
"111110001010001001010011100000000000",--981
"111110001110001001000011100000000000",--982
"111110001010000001010010100000000000",--983
"111110001010000000010010100000000000",--984
"111110001010000000110001100000000000",--985
"111110000110011000000001100000000000",--986
"111110001110001000110001100000000000",--987
"101111000001110001010011111100000000",--988
"010110001011000001100000000000000001",--989
"000100000000000000001111100000000000",--990
"111110001100010000010010100000000000",--991
"111110001100001001100011100000000000",--992
"111110001110001001000011100000000000",--993
"111110001100000001100011000000000000",--994
"111110001100000000010011000000000000",--995
"111110001100000000110001100000000000",--996
"111110000110011000000001100000000000",--997
"111110001110001000110001100000000000",--998
"101111000001110001100011111100000000",--999
"010110001101000001010000000000000001",--1000
"000100000000000000001111100000000000",--1001
"111110001010010000010011000000000000",--1002
"111110001010001001010011100000000000",--1003
"111110001110001001000011100000000000",--1004
"111110001010000001010010100000000000",--1005
"111110001010000000010010100000000000",--1006
"111110001010000000110001100000000000",--1007
"111110000110011000000001100000000000",--1008
"111110001110001000110001100000000000",--1009
"101111000001110001010011111100000000",--1010
"010110001011000001100000000000000001",--1011
"000100000000000000001111100000000000",--1012
"111110001100010000010010100000000000",--1013
"111110001100001001100011100000000000",--1014
"111110001110001001000011100000000000",--1015
"111110001100000001100011000000000000",--1016
"111110001100000000010011000000000000",--1017
"111110001100000000110001100000000000",--1018
"111110000110011000000001100000000000",--1019
"111110001110001000110001100000000000",--1020
"101110001011111000001111100000000000",--1021
"101110000111111000000010100000000000",--1022
"101110111111111000000001100000000000",--1023
"000101000000000000000000001101001100",--1024
"011011000010001111001111100000000000",--1025
"000010000000000000000001000000000000",--1026
"001001111100000000010000000000000000",--1027
"010011000101000000000000000101000101",--1028
"000010000000000000000001100000000000",--1029
"000010000000000000000010000000000000",--1030
"000010000000000000000010100000000000",--1031
"101110000001111000000001100000000000",--1032
"001001111100000000101111111111111111",--1033
"001001111100000001001111111111111110",--1034
"001001111100000000111111111111111101",--1035
"001001111100000001011111111111111100",--1036
"101001000000000000010000000000000011",--1037
"001001111100000111111111111111111011",--1038
"000111000000000000000111010110110001",--1039
"001101111100000111111111111111111011",--1040
"000011000000000000000001100000000000",--1041
"001011000010000000110000000000000000",--1042
"000011000000000000000001100000000000",--1043
"001011000010000000110000000000000001",--1044
"000011000000000000000001100000000000",--1045
"001011000010000000110000000000000010",--1046
"101110000001111000000001100000000000",--1047
"001001111100000000011111111111111011",--1048
"101001000000000000010000000000000011",--1049
"001001111100000111111111111111111010",--1050
"000111000000000000000111010110110001",--1051
"001101111100000111111111111111111010",--1052
"000011000000000000000001100000000000",--1053
"001011000010000000110000000000000000",--1054
"000011000000000000000001100000000000",--1055
"001011000010000000110000000000000001",--1056
"000011000000000000000001100000000000",--1057
"001011000010000000110000000000000010",--1058
"000011000000000000000001100000000000",--1059
"001001111100000000011111111111111010",--1060
"001011111100000000111111111111111001",--1061
"101001000000000000010000000000000010",--1062
"101110000001111000000001100000000000",--1063
"001001111100000111111111111111111000",--1064
"000111000000000000000111010110110001",--1065
"001101111100000111111111111111111000",--1066
"000011000000000000000001100000000000",--1067
"001011000010000000110000000000000000",--1068
"000011000000000000000001100000000000",--1069
"001011000010000000110000000000000001",--1070
"101110000001111000000001100000000000",--1071
"001001111100000000011111111111111000",--1072
"101001000000000000010000000000000011",--1073
"001001111100000111111111111111110111",--1074
"000111000000000000000111010110110001",--1075
"001101111100000111111111111111110111",--1076
"000011000000000000000001100000000000",--1077
"001011000010000000110000000000000000",--1078
"000011000000000000000001100000000000",--1079
"001011000010000000110000000000000001",--1080
"000011000000000000000001100000000000",--1081
"001011000010000000110000000000000010",--1082
"101110000001111000000001100000000000",--1083
"001001111100000000011111111111110111",--1084
"101001000000000000010000000000000011",--1085
"001001111100000111111111111111110110",--1086
"000111000000000000000111010110110001",--1087
"001101111100000111111111111111110110",--1088
"001101111100000000101111111111111100",--1089
"010000000101000000000000000000001111",--1090
"000011000000000000000001100000000000",--1091
"101111001001110001000011110010001110",--1092
"101111001001100001001111101000110101",--1093
"111110000110001001000001100000000000",--1094
"001011000010000000110000000000000000",--1095
"000011000000000000000001100000000000",--1096
"101111001001110001000011110010001110",--1097
"101111001001100001001111101000110101",--1098
"111110000110001001000001100000000000",--1099
"001011000010000000110000000000000001",--1100
"000011000000000000000001100000000000",--1101
"101111001001110001000011110010001110",--1102
"101111001001100001001111101000110101",--1103
"111110000110001001000001100000000000",--1104
"001011000010000000110000000000000010",--1105
"001101111100000000111111111111111101",--1106
"011111000111000000100000000000000010",--1107
"101001000000000001000000000000000001",--1108
"000101000000000000000000010001011011",--1109
"001111111100000000111111111111111001",--1110
"011010000111000000000000000000000010",--1111
"101001000000000001000000000000000001",--1112
"000101000000000000000000010001011011",--1113
"101000000001111000000010000000000000",--1114
"101110000001111000000001100000000000",--1115
"001001111100000001001111111111110110",--1116
"001001111100000000011111111111110101",--1117
"101001000000000000010000000000000100",--1118
"001001111100000111111111111111110100",--1119
"000111000000000000000111010110110001",--1120
"001101111100000111111111111111110100",--1121
"101000111011111000000001000000000000",--1122
"101001111010000111010000000000001011",--1123
"001001000100000000010000000000001010",--1124
"001101111100000000011111111111110101",--1125
"001001000100000000010000000000001001",--1126
"001101111100000000111111111111110111",--1127
"001001000100000000110000000000001000",--1128
"001101111100000000111111111111111000",--1129
"001001000100000000110000000000000111",--1130
"001101111100000000111111111111110110",--1131
"001001000100000000110000000000000110",--1132
"001101111100000000111111111111111010",--1133
"001001000100000000110000000000000101",--1134
"001101111100000000111111111111111011",--1135
"001001000100000000110000000000000100",--1136
"001101111100000001001111111111111100",--1137
"001001000100000001000000000000000011",--1138
"001101111100000001011111111111111110",--1139
"001001000100000001010000000000000010",--1140
"001101111100000001011111111111111101",--1141
"001001000100000001010000000000000001",--1142
"001101111100000001101111111111111111",--1143
"001001000100000001100000000000000000",--1144
"001101111100000001100000000000000000",--1145
"001001001100000000100000000101101101",--1146
"011111001011000000110000000000101111",--1147
"001111000110000000110000000000000000",--1148
"011110000111000000000000000000000010",--1149
"101110000001111000000001100000000000",--1150
"000101000000000000000000010010001010",--1151
"011110000111000000000000000000000010",--1152
"101110000001111000000010000000000000",--1153
"000101000000000000000000010010000111",--1154
"010110000111000000000000000000000010",--1155
"101110000011111000000010000000000000",--1156
"000101000000000000000000010010000111",--1157
"101110000101111000000010000000000000",--1158
"111110000110001000110001100000000000",--1159
"111110000110011000000001100000000000",--1160
"111110001000001000110001100000000000",--1161
"001011000110000000110000000000000000",--1162
"001111000110000000110000000000000001",--1163
"011110000111000000000000000000000010",--1164
"101110000001111000000001100000000000",--1165
"000101000000000000000000010010011001",--1166
"011110000111000000000000000000000010",--1167
"101110000001111000000010000000000000",--1168
"000101000000000000000000010010010110",--1169
"010110000111000000000000000000000010",--1170
"101110000011111000000010000000000000",--1171
"000101000000000000000000010010010110",--1172
"101110000101111000000010000000000000",--1173
"111110000110001000110001100000000000",--1174
"111110000110011000000001100000000000",--1175
"111110001000001000110001100000000000",--1176
"001011000110000000110000000000000001",--1177
"001111000110000000110000000000000010",--1178
"011110000111000000000000000000000010",--1179
"101110000001111000000001100000000000",--1180
"000101000000000000000000010010101000",--1181
"011110000111000000000000000000000010",--1182
"101110000001111000000010000000000000",--1183
"000101000000000000000000010010100101",--1184
"010110000111000000000000000000000010",--1185
"101110000011111000000010000000000000",--1186
"000101000000000000000000010010100101",--1187
"101110000101111000000010000000000000",--1188
"111110000110001000110001100000000000",--1189
"111110000110011000000001100000000000",--1190
"111110001000001000110001100000000000",--1191
"001011000110000000110000000000000010",--1192
"010000001001000000000000000010100011",--1193
"000101000000000000000000010011000111",--1194
"011111001011000000100000000000011010",--1195
"001111000110000000110000000000000000",--1196
"111110000110001000110001100000000000",--1197
"001111000110000001000000000000000001",--1198
"111110001000001001000010000000000000",--1199
"111110000110000001000001100000000000",--1200
"001111000110000001000000000000000010",--1201
"111110001000001001000010000000000000",--1202
"111110000110000001000001100000000000",--1203
"111110000110100000000001100000000000",--1204
"011110000111000000000000000000000010",--1205
"101110000011111000000001100000000000",--1206
"000101000000000000000000010010111101",--1207
"001111111100000001001111111111111001",--1208
"011010001001000000000000000000000010",--1209
"111110000110011000000001100000000000",--1210
"000101000000000000000000010010111101",--1211
"111110000110011000000001100000000010",--1212
"001111000110000001000000000000000000",--1213
"111110001000001000110010000000000000",--1214
"001011000110000001000000000000000000",--1215
"001111000110000001000000000000000001",--1216
"111110001000001000110010000000000000",--1217
"001011000110000001000000000000000001",--1218
"001111000110000001000000000000000010",--1219
"111110001000001000110001100000000000",--1220
"001011000110000000110000000000000010",--1221
"010000001001000000000000000010000110",--1222
"001111000010000000110000000000000000",--1223
"001001111100000111111111111111110100",--1224
"000111000000000000000111010110111000",--1225
"001101111100000111111111111111110100",--1226
"001101111100000000011111111111110101",--1227
"001111000010000001000000000000000000",--1228
"001011111100000000111111111111110100",--1229
"101110001001111000000001100000000000",--1230
"001001111100000111111111111111110011",--1231
"000111000000000000000111011000000010",--1232
"001101111100000111111111111111110011",--1233
"001101111100000000011111111111110101",--1234
"001111000010000001000000000000000001",--1235
"001011111100000000111111111111110011",--1236
"101110001001111000000001100000000000",--1237
"001001111100000111111111111111110010",--1238
"000111000000000000000111010110111000",--1239
"001101111100000111111111111111110010",--1240
"001101111100000000011111111111110101",--1241
"001111000010000001000000000000000001",--1242
"001011111100000000111111111111110010",--1243
"101110001001111000000001100000000000",--1244
"001001111100000111111111111111110001",--1245
"000111000000000000000111011000000010",--1246
"001101111100000111111111111111110001",--1247
"001101111100000000011111111111110101",--1248
"001111000010000001000000000000000010",--1249
"001011111100000000111111111111110001",--1250
"101110001001111000000001100000000000",--1251
"001001111100000111111111111111110000",--1252
"000111000000000000000111010110111000",--1253
"001101111100000111111111111111110000",--1254
"001101111100000000011111111111110101",--1255
"001111000010000001000000000000000010",--1256
"001011111100000000111111111111110000",--1257
"101110001001111000000001100000000000",--1258
"001001111100000111111111111111101111",--1259
"000111000000000000000111011000000010",--1260
"001101111100000111111111111111101111",--1261
"001111111100000001001111111111110000",--1262
"001111111100000001011111111111110010",--1263
"111110001010001001000011000000000000",--1264
"001111111100000001111111111111110001",--1265
"001111111100000010001111111111110011",--1266
"111110010000001001110100100000000000",--1267
"111110010010001001000100100000000000",--1268
"001111111100000010101111111111110100",--1269
"111110010100001000110101100000000000",--1270
"111110010010010010110100100000000000",--1271
"111110010100001001110101100000000000",--1272
"111110010110001001000101100000000000",--1273
"111110010000001000110110000000000000",--1274
"111110010110000011000101100000000000",--1275
"111110001010001000110110000000000000",--1276
"111110010000001001110110100000000000",--1277
"111110011010001000110110100000000000",--1278
"111110010100001001000111000000000000",--1279
"111110011010000011100110100000000000",--1280
"111110010100001001110111000000000000",--1281
"111110011100001000110001100000000000",--1282
"111110010000001001000010000000000000",--1283
"111110000110010001000001100000000000",--1284
"101110001111111000000010000000000010",--1285
"111110010000001001010011100000000000",--1286
"111110010100001001010010100000000000",--1287
"001101111100000000011111111111111011",--1288
"001111000010000010000000000000000000",--1289
"001111000010000010100000000000000001",--1290
"001111000010000011100000000000000010",--1291
"111110001100001001100111100000000000",--1292
"111110010000001011110111100000000000",--1293
"111110011000001011001000000000000000",--1294
"111110010100001100001000000000000000",--1295
"111110011110000100000111100000000000",--1296
"111110001000001001001000000000000000",--1297
"111110011100001100001000000000000000",--1298
"111110011110000100000111100000000000",--1299
"001011000010000011110000000000000000",--1300
"111110010010001010010111100000000000",--1301
"111110010000001011110111100000000000",--1302
"111110011010001011011000000000000000",--1303
"111110010100001100001000000000000000",--1304
"111110011110000100000111100000000000",--1305
"111110001110001001111000000000000000",--1306
"111110011100001100001000000000000000",--1307
"111110011110000100000111100000000000",--1308
"001011000010000011110000000000000001",--1309
"111110010110001010110111100000000000",--1310
"111110010000001011110111100000000000",--1311
"111110000110001000111000000000000000",--1312
"111110010100001100001000000000000000",--1313
"111110011110000100000111100000000000",--1314
"111110001010001001011000000000000000",--1315
"111110011100001100001000000000000000",--1316
"111110011110000100000111100000000000",--1317
"001011000010000011110000000000000010",--1318
"101111000001110011110100000000000000",--1319
"111110010000001010011000000000000000",--1320
"111110100000001010111000000000000000",--1321
"111110010100001011011000100000000000",--1322
"111110100010001000111000100000000000",--1323
"111110100000000100011000000000000000",--1324
"111110011100001001111000100000000000",--1325
"111110100010001001011000100000000000",--1326
"111110100000000100011000000000000000",--1327
"111110011110001100000111100000000000",--1328
"001101111100000000011111111111110101",--1329
"001011000010000011110000000000000000",--1330
"101111000001110011110100000000000000",--1331
"111110010000001001101000000000000000",--1332
"111110100000001010110101100000000000",--1333
"111110010100001011001000000000000000",--1334
"111110100000001000110001100000000000",--1335
"111110010110000000110001100000000000",--1336
"111110011100001001000101100000000000",--1337
"111110010110001001010010100000000000",--1338
"111110000110000001010001100000000000",--1339
"111110011110001000110001100000000000",--1340
"001011000010000000110000000000000001",--1341
"101111000001110000110100000000000000",--1342
"111110010000001001100010100000000000",--1343
"111110001010001010010010100000000000",--1344
"111110010100001011000011000000000000",--1345
"111110001100001011010011000000000000",--1346
"111110001010000001100010100000000000",--1347
"111110011100001001000010000000000000",--1348
"111110001000001001110010000000000000",--1349
"111110001010000001000010000000000000",--1350
"111110000110001001000001100000000000",--1351
"001011000010000000110000000000000010",--1352
"000101000000000000000000010101001101",--1353
"001101111100000000010000000000000000",--1354
"001001000000000000010000000110101010",--1355
"000100000000000000001111100000000000",--1356
"001101111100000000010000000000000000",--1357
"101001000010000000010000000000000001",--1358
"011011000010001111001111100000000000",--1359
"000101000000000000000000010000000010",--1360
"000010000000000000000001000000000000",--1361
"011111000101000000000000000000000011",--1362
"101001000010000000010000000000000001",--1363
"101001000000000000101111111111111111",--1364
"000101000000000000000111010110101010",--1365
"101001000010000000110000000000000001",--1366
"001001111100000000100000000000000000",--1367
"001001111100000000011111111111111111",--1368
"101000000111111000000000100000000000",--1369
"001001111100000111111111111111111110",--1370
"101001111100010111100000000000000011",--1371
"000111000000000000000000010101010001",--1372
"101001111100000111100000000000000011",--1373
"001101111100000111111111111111111110",--1374
"001101111100000000101111111111111111",--1375
"001101111100000000110000000000000000",--1376
"001000000010000000100001100000000000",--1377
"000100000000000000001111100000000000",--1378
"001001111100000000010000000000000000",--1379
"101000000001111000000000100000000000",--1380
"001001111100000111111111111111111111",--1381
"101001111100010111100000000000000010",--1382
"000111000000000000000000010101010001",--1383
"101001111100000111100000000000000010",--1384
"001101111100000111111111111111111111",--1385
"101000000011111000000001000000000000",--1386
"001101000010000000010000000000000000",--1387
"011111000011000000000000000000000011",--1388
"001101111100000000010000000000000000",--1389
"101001000010000000010000000000000001",--1390
"000101000000000000000111010110101010",--1391
"001101111100000000010000000000000000",--1392
"101001000010000000010000000000000001",--1393
"001001111100000000101111111111111111",--1394
"001001111100000111111111111111111110",--1395
"101001111100010111100000000000000011",--1396
"000111000000000000000000010101100011",--1397
"101001111100000111100000000000000011",--1398
"001101111100000111111111111111111110",--1399
"001101111100000000100000000000000000",--1400
"001101111100000000111111111111111111",--1401
"001000000010000000100001100000000000",--1402
"000100000000000000001111100000000000",--1403
"001001111100000000010000000000000000",--1404
"101000000001111000000000100000000000",--1405
"001001111100000111111111111111111111",--1406
"101001111100010111100000000000000010",--1407
"000111000000000000000000010101010001",--1408
"101001111100000111100000000000000010",--1409
"001101111100000111111111111111111111",--1410
"001101000010000000100000000000000000",--1411
"010011000100000000001111100000000000",--1412
"001101111100000000100000000000000000",--1413
"001001000100000000010000000100110001",--1414
"101001000100000000010000000000000001",--1415
"000101000000000000000000010101111100",--1416
"001101000100000000110000000101101101",--1417
"001101000010000001000000000000000001",--1418
"001101000010000001010000000000000000",--1419
"001101000110000001100000000000000001",--1420
"001001111100000000010000000000000000",--1421
"011111001101000000010000000001000111",--1422
"101110000001111000000001100000000000",--1423
"001001111100000001001111111111111111",--1424
"001001111100000000101111111111111110",--1425
"001001111100000000111111111111111101",--1426
"001001111100000001011111111111111100",--1427
"101001000000000000010000000000000110",--1428
"001001111100000111111111111111111011",--1429
"000111000000000000000111010110110001",--1430
"001101111100000111111111111111111011",--1431
"001101111100000000101111111111111100",--1432
"001111000100000000110000000000000000",--1433
"011110000111000000000000000000000010",--1434
"001011000010000000000000000000000001",--1435
"000101000000000000000000010110101100",--1436
"001101111100000000111111111111111101",--1437
"001101000110000001000000000000000110",--1438
"001111000100000000110000000000000000",--1439
"011010000111000000000000000000000010",--1440
"101001000000000001010000000000000001",--1441
"000101000000000000000000010110100100",--1442
"101000000001111000000010100000000000",--1443
"001101000110000001100000000000000100",--1444
"001111001100000000110000000000000000",--1445
"011100001001000001010000000000000001",--1446
"101110000111111000000001100000000010",--1447
"001011000010000000110000000000000000",--1448
"001111000100000000110000000000000000",--1449
"111110000110011000000001100000000000",--1450
"001011000010000000110000000000000001",--1451
"001111000100000000110000000000000001",--1452
"011110000111000000000000000000000010",--1453
"001011000010000000000000000000000011",--1454
"000101000000000000000000010110111111",--1455
"001101111100000000111111111111111101",--1456
"001101000110000001000000000000000110",--1457
"001111000100000000110000000000000001",--1458
"011010000111000000000000000000000010",--1459
"101001000000000001010000000000000001",--1460
"000101000000000000000000010110110111",--1461
"101000000001111000000010100000000000",--1462
"001101000110000001100000000000000100",--1463
"001111001100000000110000000000000001",--1464
"011100001001000001010000000000000001",--1465
"101110000111111000000001100000000010",--1466
"001011000010000000110000000000000010",--1467
"001111000100000000110000000000000001",--1468
"111110000110011000000001100000000000",--1469
"001011000010000000110000000000000011",--1470
"001111000100000000110000000000000010",--1471
"011110000111000000000000000000000010",--1472
"001011000010000000000000000000000101",--1473
"000101000000000000000000010111010010",--1474
"001101111100000000111111111111111101",--1475
"001101000110000001000000000000000110",--1476
"001111000100000000110000000000000010",--1477
"011010000111000000000000000000000010",--1478
"101001000000000001010000000000000001",--1479
"000101000000000000000000010111001010",--1480
"101000000001111000000010100000000000",--1481
"001101000110000000110000000000000100",--1482
"001111000110000000110000000000000010",--1483
"011100001001000001010000000000000001",--1484
"101110000111111000000001100000000010",--1485
"001011000010000000110000000000000100",--1486
"001111000100000000110000000000000010",--1487
"111110000110011000000001100000000000",--1488
"001011000010000000110000000000000101",--1489
"001101111100000000101111111111111110",--1490
"001101111100000001001111111111111111",--1491
"001000001000000000100000100000000000",--1492
"000101000000000000000000011001100110",--1493
"011111001101000000100000000000101100",--1494
"101110000001111000000001100000000000",--1495
"001001111100000001001111111111111111",--1496
"001001111100000000101111111111111110",--1497
"001001111100000000111111111111111101",--1498
"001001111100000001011111111111111100",--1499
"101001000000000000010000000000000100",--1500
"001001111100000111111111111111111011",--1501
"000111000000000000000111010110110001",--1502
"001101111100000111111111111111111011",--1503
"001101111100000000101111111111111100",--1504
"001111000100000000110000000000000000",--1505
"001101111100000000111111111111111101",--1506
"001101000110000000110000000000000100",--1507
"001111000110000001000000000000000000",--1508
"111110000110001001000001100000000000",--1509
"001111000100000001000000000000000001",--1510
"001111000110000001010000000000000001",--1511
"111110001000001001010010000000000000",--1512
"111110000110000001000001100000000000",--1513
"001111000100000001000000000000000010",--1514
"001111000110000001010000000000000010",--1515
"111110001000001001010010000000000000",--1516
"111110000110000001000001100000000000",--1517
"010110000111000000000000000000001111",--1518
"111110000110011000000010000000000010",--1519
"001011000010000001000000000000000000",--1520
"001111000110000001000000000000000000",--1521
"111110000110011000000010100000000000",--1522
"111110001000001001010010000000000010",--1523
"001011000010000001000000000000000001",--1524
"001111000110000001000000000000000001",--1525
"111110000110011000000010100000000000",--1526
"111110001000001001010010000000000010",--1527
"001011000010000001000000000000000010",--1528
"001111000110000001000000000000000010",--1529
"111110000110011000000001100000000000",--1530
"111110001000001000110001100000000010",--1531
"001011000010000000110000000000000011",--1532
"000101000000000000000000010111111111",--1533
"001011000010000000000000000000000000",--1534
"001101111100000000101111111111111110",--1535
"001101111100000001001111111111111111",--1536
"001000001000000000100000100000000000",--1537
"000101000000000000000000011001100110",--1538
"101110000001111000000001100000000000",--1539
"001001111100000001001111111111111111",--1540
"001001111100000000101111111111111110",--1541
"001001111100000000111111111111111101",--1542
"001001111100000001011111111111111100",--1543
"101001000000000000010000000000000101",--1544
"001001111100000111111111111111111011",--1545
"000111000000000000000111010110110001",--1546
"001101111100000111111111111111111011",--1547
"001101111100000000101111111111111100",--1548
"001111000100000000110000000000000000",--1549
"001111000100000001000000000000000001",--1550
"001111000100000001010000000000000010",--1551
"111110000110001000110011000000000000",--1552
"001101111100000000111111111111111101",--1553
"001101000110000001000000000000000100",--1554
"001111001000000001110000000000000000",--1555
"111110001100001001110011000000000000",--1556
"111110001000001001000011100000000000",--1557
"001111001000000010000000000000000001",--1558
"111110001110001010000011100000000000",--1559
"111110001100000001110011000000000000",--1560
"111110001010001001010011100000000000",--1561
"001111001000000010000000000000000010",--1562
"111110001110001010000011100000000000",--1563
"111110001100000001110011000000000000",--1564
"001101000110000001010000000000000011",--1565
"011100001011000000000000000000000010",--1566
"101110001101111000000001100000000000",--1567
"000101000000000000000000011000101110",--1568
"111110001000001001010011100000000000",--1569
"001101000110000001100000000000001001",--1570
"001111001100000010000000000000000000",--1571
"111110001110001010000011100000000000",--1572
"111110001100000001110011000000000000",--1573
"111110001010001000110010100000000000",--1574
"001111001100000001110000000000000001",--1575
"111110001010001001110010100000000000",--1576
"111110001100000001010010100000000000",--1577
"111110000110001001000001100000000000",--1578
"001111001100000001000000000000000010",--1579
"111110000110001001000001100000000000",--1580
"111110001010000000110001100000000000",--1581
"001111000100000001000000000000000000",--1582
"001111001000000001010000000000000000",--1583
"111110001000001001010010000000000010",--1584
"001111000100000001010000000000000001",--1585
"001111001000000001100000000000000001",--1586
"111110001010001001100010100000000010",--1587
"001111000100000001100000000000000010",--1588
"001111001000000001110000000000000010",--1589
"111110001100001001110011000000000010",--1590
"001011000010000000110000000000000000",--1591
"011100001011000000000000000000000101",--1592
"001011000010000001000000000000000001",--1593
"001011000010000001010000000000000010",--1594
"001011000010000001100000000000000011",--1595
"010010000111000000000000000000100110",--1596
"000101000000000000000000011001100001",--1597
"001111000100000001110000000000000010",--1598
"001101000110000000110000000000001001",--1599
"001111000110000010000000000000000001",--1600
"111110001110001010000011100000000000",--1601
"001111000100000010000000000000000001",--1602
"001111000110000010010000000000000010",--1603
"111110010000001010010100000000000000",--1604
"111110001110000010000011100000000000",--1605
"101111000001110010000011111100000000",--1606
"111110001110001010000011100000000000",--1607
"111110001000010001110010000000000000",--1608
"001011000010000001000000000000000001",--1609
"001111000100000001000000000000000010",--1610
"001111000110000001110000000000000000",--1611
"111110001000001001110010000000000000",--1612
"001111000100000001110000000000000000",--1613
"001111000110000010000000000000000010",--1614
"111110001110001010000011100000000000",--1615
"111110001000000001110010000000000000",--1616
"101111000001110001110011111100000000",--1617
"111110001000001001110010000000000000",--1618
"111110001010010001000010000000000000",--1619
"001011000010000001000000000000000010",--1620
"001111000100000001000000000000000001",--1621
"001111000110000001010000000000000000",--1622
"111110001000001001010010000000000000",--1623
"001111000100000001010000000000000000",--1624
"001111000110000001110000000000000001",--1625
"111110001010001001110010100000000000",--1626
"111110001000000001010010000000000000",--1627
"101111000001110001010011111100000000",--1628
"111110001000001001010010000000000000",--1629
"111110001100010001000010000000000000",--1630
"001011000010000001000000000000000011",--1631
"010010000111000000000000000000000010",--1632
"111110000110011000000001100000000000",--1633
"001011000010000000110000000000000100",--1634
"001101111100000000101111111111111110",--1635
"001101111100000001001111111111111111",--1636
"001000001000000000100000100000000000",--1637
"101001000100010000100000000000000001",--1638
"001101111100000000010000000000000000",--1639
"010111000100000000001111100000000000",--1640
"000101000000000000000000010110001001",--1641
"001101000000000000100000000110101010",--1642
"101001000100010000100000000000000001",--1643
"010111000100000000001111100000000000",--1644
"000101000000000000000000010110001001",--1645
"010111000100000000001111100000000000",--1646
"001101000100000000110000000101101101",--1647
"001101000110000001000000000000001010",--1648
"001101000110000001010000000000000001",--1649
"001111000010000000110000000000000000",--1650
"001101000110000001100000000000000101",--1651
"001111001100000001000000000000000000",--1652
"111110000110010001000001100000000000",--1653
"001011001000000000110000000000000000",--1654
"001111000010000000110000000000000001",--1655
"001111001100000001000000000000000001",--1656
"111110000110010001000001100000000000",--1657
"001011001000000000110000000000000001",--1658
"001111000010000000110000000000000010",--1659
"001111001100000001000000000000000010",--1660
"111110000110010001000001100000000000",--1661
"001011001000000000110000000000000010",--1662
"011111001011000000100000000000001110",--1663
"001101000110000000110000000000000100",--1664
"001111001000000000110000000000000000",--1665
"001111001000000001000000000000000001",--1666
"001111001000000001010000000000000010",--1667
"001111000110000001100000000000000000",--1668
"111110001100001000110001100000000000",--1669
"001111000110000001100000000000000001",--1670
"111110001100001001000010000000000000",--1671
"111110000110000001000001100000000000",--1672
"001111000110000001000000000000000010",--1673
"111110001000001001010010000000000000",--1674
"111110000110000001000001100000000000",--1675
"001011001000000000110000000000000011",--1676
"000101000000000000000000011010110011",--1677
"010111001011000000100000000000100100",--1678
"001111001000000000110000000000000000",--1679
"001111001000000001000000000000000001",--1680
"001111001000000001010000000000000010",--1681
"111110000110001000110011000000000000",--1682
"001101000110000001100000000000000100",--1683
"001111001100000001110000000000000000",--1684
"111110001100001001110011000000000000",--1685
"111110001000001001000011100000000000",--1686
"001111001100000010000000000000000001",--1687
"111110001110001010000011100000000000",--1688
"111110001100000001110011000000000000",--1689
"111110001010001001010011100000000000",--1690
"001111001100000010000000000000000010",--1691
"111110001110001010000011100000000000",--1692
"111110001100000001110011000000000000",--1693
"001101000110000001100000000000000011",--1694
"011100001101000000000000000000000011",--1695
"101110001101111000000001100000000000",--1696
"011111001011000000110000000000010000",--1697
"000101000000000000000000011010110001",--1698
"111110001000001001010011100000000000",--1699
"001101000110000000110000000000001001",--1700
"001111000110000010000000000000000000",--1701
"111110001110001010000011100000000000",--1702
"111110001100000001110011000000000000",--1703
"111110001010001000110010100000000000",--1704
"001111000110000001110000000000000001",--1705
"111110001010001001110010100000000000",--1706
"111110001100000001010010100000000000",--1707
"111110000110001001000001100000000000",--1708
"001111000110000001000000000000000010",--1709
"111110000110001001000001100000000000",--1710
"111110001010000000110001100000000000",--1711
"011111001011000000110000000000000001",--1712
"111110000110010000010001100000000000",--1713
"001011001000000000110000000000000011",--1714
"101001000100010000100000000000000001",--1715
"010111000100000000001111100000000000",--1716
"001101000100000000110000000101101101",--1717
"001101000110000001000000000000001010",--1718
"001101000110000001010000000000000001",--1719
"001111000010000000110000000000000000",--1720
"001101000110000001100000000000000101",--1721
"001111001100000001000000000000000000",--1722
"111110000110010001000001100000000000",--1723
"001011001000000000110000000000000000",--1724
"001111000010000000110000000000000001",--1725
"001111001100000001000000000000000001",--1726
"111110000110010001000001100000000000",--1727
"001011001000000000110000000000000001",--1728
"001111000010000000110000000000000010",--1729
"001111001100000001000000000000000010",--1730
"111110000110010001000001100000000000",--1731
"001011001000000000110000000000000010",--1732
"011111001011000000100000000000001110",--1733
"001101000110000000110000000000000100",--1734
"001111001000000000110000000000000000",--1735
"001111001000000001000000000000000001",--1736
"001111001000000001010000000000000010",--1737
"001111000110000001100000000000000000",--1738
"111110001100001000110001100000000000",--1739
"001111000110000001100000000000000001",--1740
"111110001100001001000010000000000000",--1741
"111110000110000001000001100000000000",--1742
"001111000110000001000000000000000010",--1743
"111110001000001001010010000000000000",--1744
"111110000110000001000001100000000000",--1745
"001011001000000000110000000000000011",--1746
"000101000000000000000000011011111001",--1747
"010111001011000000100000000000100100",--1748
"001111001000000000110000000000000000",--1749
"001111001000000001000000000000000001",--1750
"001111001000000001010000000000000010",--1751
"111110000110001000110011000000000000",--1752
"001101000110000001100000000000000100",--1753
"001111001100000001110000000000000000",--1754
"111110001100001001110011000000000000",--1755
"111110001000001001000011100000000000",--1756
"001111001100000010000000000000000001",--1757
"111110001110001010000011100000000000",--1758
"111110001100000001110011000000000000",--1759
"111110001010001001010011100000000000",--1760
"001111001100000010000000000000000010",--1761
"111110001110001010000011100000000000",--1762
"111110001100000001110011000000000000",--1763
"001101000110000001100000000000000011",--1764
"011100001101000000000000000000000011",--1765
"101110001101111000000001100000000000",--1766
"011111001011000000110000000000010000",--1767
"000101000000000000000000011011110111",--1768
"111110001000001001010011100000000000",--1769
"001101000110000000110000000000001001",--1770
"001111000110000010000000000000000000",--1771
"111110001110001010000011100000000000",--1772
"111110001100000001110011000000000000",--1773
"111110001010001000110010100000000000",--1774
"001111000110000001110000000000000001",--1775
"111110001010001001110010100000000000",--1776
"111110001100000001010010100000000000",--1777
"111110000110001001000001100000000000",--1778
"001111000110000001000000000000000010",--1779
"111110000110001001000001100000000000",--1780
"111110001010000000110001100000000000",--1781
"011111001011000000110000000000000001",--1782
"111110000110010000010001100000000000",--1783
"001011001000000000110000000000000011",--1784
"101001000100010000100000000000000001",--1785
"010111000100000000001111100000000000",--1786
"001101000100000000110000000101101101",--1787
"001101000110000001000000000000001010",--1788
"001101000110000001010000000000000001",--1789
"001111000010000000110000000000000000",--1790
"001101000110000001100000000000000101",--1791
"001111001100000001000000000000000000",--1792
"111110000110010001000001100000000000",--1793
"001011001000000000110000000000000000",--1794
"001111000010000000110000000000000001",--1795
"001111001100000001000000000000000001",--1796
"111110000110010001000001100000000000",--1797
"001011001000000000110000000000000001",--1798
"001111000010000000110000000000000010",--1799
"001111001100000001000000000000000010",--1800
"111110000110010001000001100000000000",--1801
"001011001000000000110000000000000010",--1802
"011111001011000000100000000000001110",--1803
"001101000110000000110000000000000100",--1804
"001111001000000000110000000000000000",--1805
"001111001000000001000000000000000001",--1806
"001111001000000001010000000000000010",--1807
"001111000110000001100000000000000000",--1808
"111110001100001000110001100000000000",--1809
"001111000110000001100000000000000001",--1810
"111110001100001001000010000000000000",--1811
"111110000110000001000001100000000000",--1812
"001111000110000001000000000000000010",--1813
"111110001000001001010010000000000000",--1814
"111110000110000001000001100000000000",--1815
"001011001000000000110000000000000011",--1816
"000101000000000000000000011100111111",--1817
"010111001011000000100000000000100100",--1818
"001111001000000000110000000000000000",--1819
"001111001000000001000000000000000001",--1820
"001111001000000001010000000000000010",--1821
"111110000110001000110011000000000000",--1822
"001101000110000001100000000000000100",--1823
"001111001100000001110000000000000000",--1824
"111110001100001001110011000000000000",--1825
"111110001000001001000011100000000000",--1826
"001111001100000010000000000000000001",--1827
"111110001110001010000011100000000000",--1828
"111110001100000001110011000000000000",--1829
"111110001010001001010011100000000000",--1830
"001111001100000010000000000000000010",--1831
"111110001110001010000011100000000000",--1832
"111110001100000001110011000000000000",--1833
"001101000110000001100000000000000011",--1834
"011100001101000000000000000000000011",--1835
"101110001101111000000001100000000000",--1836
"011111001011000000110000000000010000",--1837
"000101000000000000000000011100111101",--1838
"111110001000001001010011100000000000",--1839
"001101000110000000110000000000001001",--1840
"001111000110000010000000000000000000",--1841
"111110001110001010000011100000000000",--1842
"111110001100000001110011000000000000",--1843
"111110001010001000110010100000000000",--1844
"001111000110000001110000000000000001",--1845
"111110001010001001110010100000000000",--1846
"111110001100000001010010100000000000",--1847
"111110000110001001000001100000000000",--1848
"001111000110000001000000000000000010",--1849
"111110000110001001000001100000000000",--1850
"111110001010000000110001100000000000",--1851
"011111001011000000110000000000000001",--1852
"111110000110010000010001100000000000",--1853
"001011001000000000110000000000000011",--1854
"101001000100010000100000000000000001",--1855
"010111000100000000001111100000000000",--1856
"001101000100000000110000000101101101",--1857
"001101000110000001000000000000001010",--1858
"001101000110000001010000000000000001",--1859
"001111000010000000110000000000000000",--1860
"001101000110000001100000000000000101",--1861
"001111001100000001000000000000000000",--1862
"111110000110010001000001100000000000",--1863
"001011001000000000110000000000000000",--1864
"001111000010000000110000000000000001",--1865
"001111001100000001000000000000000001",--1866
"111110000110010001000001100000000000",--1867
"001011001000000000110000000000000001",--1868
"001111000010000000110000000000000010",--1869
"001111001100000001000000000000000010",--1870
"111110000110010001000001100000000000",--1871
"001011001000000000110000000000000010",--1872
"011111001011000000100000000000001110",--1873
"001101000110000000110000000000000100",--1874
"001111001000000000110000000000000000",--1875
"001111001000000001000000000000000001",--1876
"001111001000000001010000000000000010",--1877
"001111000110000001100000000000000000",--1878
"111110001100001000110001100000000000",--1879
"001111000110000001100000000000000001",--1880
"111110001100001001000010000000000000",--1881
"111110000110000001000001100000000000",--1882
"001111000110000001000000000000000010",--1883
"111110001000001001010010000000000000",--1884
"111110000110000001000001100000000000",--1885
"001011001000000000110000000000000011",--1886
"000101000000000000000000011110000101",--1887
"010111001011000000100000000000100100",--1888
"001111001000000000110000000000000000",--1889
"001111001000000001000000000000000001",--1890
"001111001000000001010000000000000010",--1891
"111110000110001000110011000000000000",--1892
"001101000110000001100000000000000100",--1893
"001111001100000001110000000000000000",--1894
"111110001100001001110011000000000000",--1895
"111110001000001001000011100000000000",--1896
"001111001100000010000000000000000001",--1897
"111110001110001010000011100000000000",--1898
"111110001100000001110011000000000000",--1899
"111110001010001001010011100000000000",--1900
"001111001100000010000000000000000010",--1901
"111110001110001010000011100000000000",--1902
"111110001100000001110011000000000000",--1903
"001101000110000001100000000000000011",--1904
"011100001101000000000000000000000011",--1905
"101110001101111000000001100000000000",--1906
"011111001011000000110000000000010000",--1907
"000101000000000000000000011110000011",--1908
"111110001000001001010011100000000000",--1909
"001101000110000000110000000000001001",--1910
"001111000110000010000000000000000000",--1911
"111110001110001010000011100000000000",--1912
"111110001100000001110011000000000000",--1913
"111110001010001000110010100000000000",--1914
"001111000110000001110000000000000001",--1915
"111110001010001001110010100000000000",--1916
"111110001100000001010010100000000000",--1917
"111110000110001001000001100000000000",--1918
"001111000110000001000000000000000010",--1919
"111110000110001001000001100000000000",--1920
"111110001010000000110001100000000000",--1921
"011111001011000000110000000000000001",--1922
"111110000110010000010001100000000000",--1923
"001011001000000000110000000000000011",--1924
"101001000100010000100000000000000001",--1925
"010111000100000000001111100000000000",--1926
"000101000000000000000000011001101111",--1927
"001100000100000000010001100000000000",--1928
"011111000111000000000000000000000010",--1929
"101001000000000000010000000000000001",--1930
"000100000000000000001111100000000000",--1931
"001101000110000000110000000101101101",--1932
"001101000110000001000000000000000101",--1933
"001111001000000001100000000000000000",--1934
"111110000110010001100011000000000000",--1935
"001111001000000001110000000000000001",--1936
"111110001000010001110011100000000000",--1937
"001111001000000010000000000000000010",--1938
"111110001010010010000100000000000000",--1939
"001101000110000001000000000000000001",--1940
"011111001001000000010000000000010000",--1941
"101110001101111000000011000000000001",--1942
"001101000110000001000000000000000100",--1943
"001111001000000010010000000000000000",--1944
"010110010011000001100000000000001001",--1945
"101110001111111000000011000000000001",--1946
"001111001000000001110000000000000001",--1947
"010110001111000001100000000000000110",--1948
"101110010001111000000011000000000001",--1949
"001111001000000001110000000000000010",--1950
"010110001111000001100000000000000011",--1951
"001101000110000000110000000000000110",--1952
"011100000111000000000000000100111101",--1953
"000101000000000000000000011111011011",--1954
"001101000110000000110000000000000110",--1955
"011100000111000000000000000000110110",--1956
"000101000000000000000000100011011111",--1957
"011111001001000000100000000000001111",--1958
"001101000110000001000000000000000100",--1959
"001111001000000010010000000000000000",--1960
"111110010010001001100011000000000000",--1961
"001111001000000010010000000000000001",--1962
"111110010010001001110011100000000000",--1963
"111110001100000001110011000000000000",--1964
"001111001000000001110000000000000010",--1965
"111110001110001010000011100000000000",--1966
"111110001100000001110011000000000000",--1967
"001101000110000000110000000000000110",--1968
"011010001101000000000000000000000010",--1969
"011111000111000000010000000000101000",--1970
"000101000000000000000000100011011111",--1971
"011100000111000000000000000000100110",--1972
"000101000000000000000000100011011111",--1973
"111110001100001001100100100000000000",--1974
"001101000110000001010000000000000100",--1975
"001111001010000010100000000000000000",--1976
"111110010010001010100100100000000000",--1977
"111110001110001001110101000000000000",--1978
"001111001010000010110000000000000001",--1979
"111110010100001010110101000000000000",--1980
"111110010010000010100100100000000000",--1981
"111110010000001010000101000000000000",--1982
"001111001010000010110000000000000010",--1983
"111110010100001010110101000000000000",--1984
"111110010010000010100100100000000000",--1985
"001101000110000001010000000000000011",--1986
"011100001011000000000000000000000011",--1987
"101110010011111000000011000000000000",--1988
"011111001001000000110000000000010000",--1989
"000101000000000000000000011111010101",--1990
"111110001110001010000101000000000000",--1991
"001101000110000001010000000000001001",--1992
"001111001010000010110000000000000000",--1993
"111110010100001010110101000000000000",--1994
"111110010010000010100100100000000000",--1995
"111110010000001001100100000000000000",--1996
"001111001010000010100000000000000001",--1997
"111110010000001010100100000000000000",--1998
"111110010010000010000100000000000000",--1999
"111110001100001001110011000000000000",--2000
"001111001010000001110000000000000010",--2001
"111110001100001001110011000000000000",--2002
"111110010000000001100011000000000000",--2003
"011111001001000000110000000000000001",--2004
"111110001100010000010011000000000000",--2005
"001101000110000000110000000000000110",--2006
"011010001101000000000000000000000010",--2007
"011111000111000000010000000000000010",--2008
"000101000000000000000000100011011111",--2009
"010000000111000000000000000100000100",--2010
"101001000010000000010000000000000001",--2011
"001100000100000000010001100000000000",--2012
"011111000111000000000000000000000010",--2013
"101001000000000000010000000000000001",--2014
"000100000000000000001111100000000000",--2015
"001101000110000000110000000101101101",--2016
"001101000110000001000000000000000101",--2017
"001111001000000001100000000000000000",--2018
"111110000110010001100011000000000000",--2019
"001111001000000001110000000000000001",--2020
"111110001000010001110011100000000000",--2021
"001111001000000010000000000000000010",--2022
"111110001010010010000100000000000000",--2023
"001101000110000001000000000000000001",--2024
"011111001001000000010000000000010000",--2025
"101110001101111000000011000000000001",--2026
"001101000110000001000000000000000100",--2027
"001111001000000010010000000000000000",--2028
"010110010011000001100000000000001001",--2029
"101110001111111000000011000000000001",--2030
"001111001000000001110000000000000001",--2031
"010110001111000001100000000000000110",--2032
"101110010001111000000011000000000001",--2033
"001111001000000001110000000000000010",--2034
"010110001111000001100000000000000011",--2035
"001101000110000000110000000000000110",--2036
"011100000111000000000000000011100111",--2037
"000101000000000000000000100000101111",--2038
"001101000110000000110000000000000110",--2039
"011100000111000000000000000000110110",--2040
"000101000000000000000000100011011101",--2041
"011111001001000000100000000000001111",--2042
"001101000110000001000000000000000100",--2043
"001111001000000010010000000000000000",--2044
"111110010010001001100011000000000000",--2045
"001111001000000010010000000000000001",--2046
"111110010010001001110011100000000000",--2047
"111110001100000001110011000000000000",--2048
"001111001000000001110000000000000010",--2049
"111110001110001010000011100000000000",--2050
"111110001100000001110011000000000000",--2051
"001101000110000000110000000000000110",--2052
"011010001101000000000000000000000010",--2053
"011111000111000000010000000000101000",--2054
"000101000000000000000000100011011101",--2055
"011100000111000000000000000000100110",--2056
"000101000000000000000000100011011101",--2057
"111110001100001001100100100000000000",--2058
"001101000110000001010000000000000100",--2059
"001111001010000010100000000000000000",--2060
"111110010010001010100100100000000000",--2061
"111110001110001001110101000000000000",--2062
"001111001010000010110000000000000001",--2063
"111110010100001010110101000000000000",--2064
"111110010010000010100100100000000000",--2065
"111110010000001010000101000000000000",--2066
"001111001010000010110000000000000010",--2067
"111110010100001010110101000000000000",--2068
"111110010010000010100100100000000000",--2069
"001101000110000001010000000000000011",--2070
"011100001011000000000000000000000011",--2071
"101110010011111000000011000000000000",--2072
"011111001001000000110000000000010000",--2073
"000101000000000000000000100000101001",--2074
"111110001110001010000101000000000000",--2075
"001101000110000001010000000000001001",--2076
"001111001010000010110000000000000000",--2077
"111110010100001010110101000000000000",--2078
"111110010010000010100100100000000000",--2079
"111110010000001001100100000000000000",--2080
"001111001010000010100000000000000001",--2081
"111110010000001010100100000000000000",--2082
"111110010010000010000100000000000000",--2083
"111110001100001001110011000000000000",--2084
"001111001010000001110000000000000010",--2085
"111110001100001001110011000000000000",--2086
"111110010000000001100011000000000000",--2087
"011111001001000000110000000000000001",--2088
"111110001100010000010011000000000000",--2089
"001101000110000000110000000000000110",--2090
"011010001101000000000000000000000010",--2091
"011111000111000000010000000000000010",--2092
"000101000000000000000000100011011101",--2093
"010000000111000000000000000010101110",--2094
"101001000010000000010000000000000001",--2095
"001100000100000000010001100000000000",--2096
"011111000111000000000000000000000010",--2097
"101001000000000000010000000000000001",--2098
"000100000000000000001111100000000000",--2099
"001101000110000000110000000101101101",--2100
"001101000110000001000000000000000101",--2101
"001111001000000001100000000000000000",--2102
"111110000110010001100011000000000000",--2103
"001111001000000001110000000000000001",--2104
"111110001000010001110011100000000000",--2105
"001111001000000010000000000000000010",--2106
"111110001010010010000100000000000000",--2107
"001101000110000001000000000000000001",--2108
"011111001001000000010000000000010000",--2109
"101110001101111000000011000000000001",--2110
"001101000110000001000000000000000100",--2111
"001111001000000010010000000000000000",--2112
"010110010011000001100000000000001001",--2113
"101110001111111000000011000000000001",--2114
"001111001000000001110000000000000001",--2115
"010110001111000001100000000000000110",--2116
"101110010001111000000011000000000001",--2117
"001111001000000001110000000000000010",--2118
"010110001111000001100000000000000011",--2119
"001101000110000000110000000000000110",--2120
"011100000111000000000000000010010001",--2121
"000101000000000000000000100010000011",--2122
"001101000110000000110000000000000110",--2123
"011100000111000000000000000000110110",--2124
"000101000000000000000000100011011011",--2125
"011111001001000000100000000000001111",--2126
"001101000110000001000000000000000100",--2127
"001111001000000010010000000000000000",--2128
"111110010010001001100011000000000000",--2129
"001111001000000010010000000000000001",--2130
"111110010010001001110011100000000000",--2131
"111110001100000001110011000000000000",--2132
"001111001000000001110000000000000010",--2133
"111110001110001010000011100000000000",--2134
"111110001100000001110011000000000000",--2135
"001101000110000000110000000000000110",--2136
"011010001101000000000000000000000010",--2137
"011111000111000000010000000000101000",--2138
"000101000000000000000000100011011011",--2139
"011100000111000000000000000000100110",--2140
"000101000000000000000000100011011011",--2141
"111110001100001001100100100000000000",--2142
"001101000110000001010000000000000100",--2143
"001111001010000010100000000000000000",--2144
"111110010010001010100100100000000000",--2145
"111110001110001001110101000000000000",--2146
"001111001010000010110000000000000001",--2147
"111110010100001010110101000000000000",--2148
"111110010010000010100100100000000000",--2149
"111110010000001010000101000000000000",--2150
"001111001010000010110000000000000010",--2151
"111110010100001010110101000000000000",--2152
"111110010010000010100100100000000000",--2153
"001101000110000001010000000000000011",--2154
"011100001011000000000000000000000011",--2155
"101110010011111000000011000000000000",--2156
"011111001001000000110000000000010000",--2157
"000101000000000000000000100001111101",--2158
"111110001110001010000101000000000000",--2159
"001101000110000001010000000000001001",--2160
"001111001010000010110000000000000000",--2161
"111110010100001010110101000000000000",--2162
"111110010010000010100100100000000000",--2163
"111110010000001001100100000000000000",--2164
"001111001010000010100000000000000001",--2165
"111110010000001010100100000000000000",--2166
"111110010010000010000100000000000000",--2167
"111110001100001001110011000000000000",--2168
"001111001010000001110000000000000010",--2169
"111110001100001001110011000000000000",--2170
"111110010000000001100011000000000000",--2171
"011111001001000000110000000000000001",--2172
"111110001100010000010011000000000000",--2173
"001101000110000000110000000000000110",--2174
"011010001101000000000000000000000010",--2175
"011111000111000000010000000000000010",--2176
"000101000000000000000000100011011011",--2177
"010000000111000000000000000001011000",--2178
"101001000010000000010000000000000001",--2179
"001100000100000000010001100000000000",--2180
"011111000111000000000000000000000010",--2181
"101001000000000000010000000000000001",--2182
"000100000000000000001111100000000000",--2183
"001101000110000000110000000101101101",--2184
"001101000110000001000000000000000101",--2185
"001111001000000001100000000000000000",--2186
"111110000110010001100011000000000000",--2187
"001111001000000001110000000000000001",--2188
"111110001000010001110011100000000000",--2189
"001111001000000010000000000000000010",--2190
"111110001010010010000100000000000000",--2191
"001101000110000001000000000000000001",--2192
"011111001001000000010000000000010000",--2193
"101110001101111000000011000000000001",--2194
"001101000110000001000000000000000100",--2195
"001111001000000010010000000000000000",--2196
"010110010011000001100000000000001001",--2197
"101110001111111000000011000000000001",--2198
"001111001000000001110000000000000001",--2199
"010110001111000001100000000000000110",--2200
"101110010001111000000011000000000001",--2201
"001111001000000001110000000000000010",--2202
"010110001111000001100000000000000011",--2203
"001101000110000000110000000000000110",--2204
"011100000111000000000000000000111011",--2205
"000101000000000000000000100011010111",--2206
"001101000110000000110000000000000110",--2207
"011100000111000000000000000000110110",--2208
"000101000000000000000000100011011001",--2209
"011111001001000000100000000000001111",--2210
"001101000110000001000000000000000100",--2211
"001111001000000010010000000000000000",--2212
"111110010010001001100011000000000000",--2213
"001111001000000010010000000000000001",--2214
"111110010010001001110011100000000000",--2215
"111110001100000001110011000000000000",--2216
"001111001000000001110000000000000010",--2217
"111110001110001010000011100000000000",--2218
"111110001100000001110011000000000000",--2219
"001101000110000000110000000000000110",--2220
"011010001101000000000000000000000010",--2221
"011111000111000000010000000000101000",--2222
"000101000000000000000000100011011001",--2223
"011100000111000000000000000000100110",--2224
"000101000000000000000000100011011001",--2225
"111110001100001001100100100000000000",--2226
"001101000110000001010000000000000100",--2227
"001111001010000010100000000000000000",--2228
"111110010010001010100100100000000000",--2229
"111110001110001001110101000000000000",--2230
"001111001010000010110000000000000001",--2231
"111110010100001010110101000000000000",--2232
"111110010010000010100100100000000000",--2233
"111110010000001010000101000000000000",--2234
"001111001010000010110000000000000010",--2235
"111110010100001010110101000000000000",--2236
"111110010010000010100100100000000000",--2237
"001101000110000001010000000000000011",--2238
"011100001011000000000000000000000011",--2239
"101110010011111000000011000000000000",--2240
"011111001001000000110000000000010000",--2241
"000101000000000000000000100011010001",--2242
"111110001110001010000101000000000000",--2243
"001101000110000001010000000000001001",--2244
"001111001010000010110000000000000000",--2245
"111110010100001010110101000000000000",--2246
"111110010010000010100100100000000000",--2247
"111110010000001001100100000000000000",--2248
"001111001010000010100000000000000001",--2249
"111110010000001010100100000000000000",--2250
"111110010010000010000100000000000000",--2251
"111110001100001001110011000000000000",--2252
"001111001010000001110000000000000010",--2253
"111110001100001001110011000000000000",--2254
"111110010000000001100011000000000000",--2255
"011111001001000000110000000000000001",--2256
"111110001100010000010011000000000000",--2257
"001101000110000000110000000000000110",--2258
"011010001101000000000000000000000010",--2259
"011111000111000000010000000000000010",--2260
"000101000000000000000000100011011001",--2261
"010000000111000000000000000000000010",--2262
"101001000010000000010000000000000001",--2263
"000101000000000000000000011110001000",--2264
"101000000001111000000000100000000000",--2265
"000100000000000000001111100000000000",--2266
"101000000001111000000000100000000000",--2267
"000100000000000000001111100000000000",--2268
"101000000001111000000000100000000000",--2269
"000100000000000000001111100000000000",--2270
"101000000001111000000000100000000000",--2271
"000100000000000000001111100000000000",--2272
"001100000100000000010001100000000000",--2273
"011111000111000000000000000000000010",--2274
"101000000001111000000000100000000000",--2275
"000100000000000000001111100000000000",--2276
"001100000100000000010001100000000000",--2277
"001101000110000001000000000101101101",--2278
"001111000000000000110000000100101010",--2279
"001101001000000001010000000000000101",--2280
"001111001010000001000000000000000000",--2281
"111110000110010001000001100000000000",--2282
"001111000000000001000000000100101011",--2283
"001111001010000001010000000000000001",--2284
"111110001000010001010010000000000000",--2285
"001111000000000001010000000100101100",--2286
"001111001010000001100000000000000010",--2287
"111110001010010001100010100000000000",--2288
"001101000110000001010000000010111110",--2289
"001101001000000001100000000000000001",--2290
"011111001101000000010000000000111100",--2291
"001111001010000001100000000000000000",--2292
"111110001100010000110011000000000000",--2293
"001111001010000001110000000000000001",--2294
"111110001100001001110011000000000000",--2295
"001111000000000001110000000011111011",--2296
"111110001100001001110011100000000000",--2297
"111110001110000001000011100000000001",--2298
"001101001000000001000000000000000100",--2299
"001111001000000010000000000000000001",--2300
"010110010001000001110000000000000111",--2301
"001111000000000001110000000011111100",--2302
"111110001100001001110011100000000000",--2303
"111110001110000001010011100000000001",--2304
"001111001000000010000000000000000010",--2305
"010110010001000001110000000000000010",--2306
"001111001010000001110000000000000001",--2307
"011110001111000000000000000000101000",--2308
"001111001010000001100000000000000010",--2309
"111110001100010001000011000000000000",--2310
"001111001010000001110000000000000011",--2311
"111110001100001001110011000000000000",--2312
"001111000000000001110000000011111010",--2313
"111110001100001001110011100000000000",--2314
"111110001110000000110011100000000001",--2315
"001111001000000010000000000000000000",--2316
"010110010001000001110000000000000111",--2317
"001111000000000001110000000011111100",--2318
"111110001100001001110011100000000000",--2319
"111110001110000001010011100000000001",--2320
"001111001000000010000000000000000010",--2321
"010110010001000001110000000000000010",--2322
"001111001010000001110000000000000011",--2323
"011110001111000000000000000000010101",--2324
"001111001010000001100000000000000100",--2325
"111110001100010001010010100000000000",--2326
"001111001010000001100000000000000101",--2327
"111110001010001001100010100000000000",--2328
"001111000000000001100000000011111010",--2329
"111110001010001001100011000000000000",--2330
"111110001100000000110001100000000001",--2331
"001111001000000001100000000000000000",--2332
"010110001101000000110000000000000111",--2333
"001111000000000000110000000011111011",--2334
"111110001010001000110001100000000000",--2335
"111110000110000001000001100000000001",--2336
"001111001000000001000000000000000001",--2337
"010110001001000000110000000000000010",--2338
"001111001010000000110000000000000101",--2339
"011110000111000000000000000000000010",--2340
"101000000001111000000010000000000000",--2341
"000101000000000000000000100110000000",--2342
"001011000000000001010000000100101111",--2343
"101001000000000001000000000000000011",--2344
"000101000000000000000000100110000000",--2345
"001011000000000001100000000100101111",--2346
"101001000000000001000000000000000010",--2347
"000101000000000000000000100110000000",--2348
"001011000000000001100000000100101111",--2349
"101001000000000001000000000000000001",--2350
"000101000000000000000000100110000000",--2351
"011111001101000000100000000000001111",--2352
"001111001010000001100000000000000000",--2353
"011010001101000000000000000000001011",--2354
"001111001010000001100000000000000001",--2355
"111110001100001000110001100000000000",--2356
"001111001010000001100000000000000010",--2357
"111110001100001001000010000000000000",--2358
"111110000110000001000001100000000000",--2359
"001111001010000001000000000000000011",--2360
"111110001000001001010010000000000000",--2361
"111110000110000001000001100000000000",--2362
"001011000000000000110000000100101111",--2363
"101001000000000001000000000000000001",--2364
"000101000000000000000000100110000000",--2365
"101000000001111000000010000000000000",--2366
"000101000000000000000000100110000000",--2367
"001111001010000001100000000000000000",--2368
"011110001101000000000000000000000010",--2369
"101000000001111000000010000000000000",--2370
"000101000000000000000000100110000000",--2371
"001111001010000001110000000000000001",--2372
"111110001110001000110011100000000000",--2373
"001111001010000010000000000000000010",--2374
"111110010000001001000100000000000000",--2375
"111110001110000010000011100000000000",--2376
"001111001010000010000000000000000011",--2377
"111110010000001001010100000000000000",--2378
"111110001110000010000011100000000000",--2379
"111110000110001000110100000000000000",--2380
"001101001000000001110000000000000100",--2381
"001111001110000010010000000000000000",--2382
"111110010000001010010100000000000000",--2383
"111110001000001001000100100000000000",--2384
"001111001110000010100000000000000001",--2385
"111110010010001010100100100000000000",--2386
"111110010000000010010100000000000000",--2387
"111110001010001001010100100000000000",--2388
"001111001110000010100000000000000010",--2389
"111110010010001010100100100000000000",--2390
"111110010000000010010100000000000000",--2391
"001101001000000001110000000000000011",--2392
"011100001111000000000000000000000011",--2393
"101110010001111000000001100000000000",--2394
"011111001101000000110000000000010000",--2395
"000101000000000000000000100101101011",--2396
"111110001000001001010100100000000000",--2397
"001101001000000001110000000000001001",--2398
"001111001110000010100000000000000000",--2399
"111110010010001010100100100000000000",--2400
"111110010000000010010100000000000000",--2401
"111110001010001000110010100000000000",--2402
"001111001110000010010000000000000001",--2403
"111110001010001010010010100000000000",--2404
"111110010000000001010010100000000000",--2405
"111110000110001001000001100000000000",--2406
"001111001110000001000000000000000010",--2407
"111110000110001001000001100000000000",--2408
"111110001010000000110001100000000000",--2409
"011111001101000000110000000000000001",--2410
"111110000110010000010001100000000000",--2411
"111110001110001001110010000000000000",--2412
"111110001100001000110001100000000000",--2413
"111110001000010000110001100000000000",--2414
"010110000111000000000000000000001111",--2415
"001101001000000001000000000000000110",--2416
"011100001001000000000000000000000110",--2417
"111110000110100000000001100000000000",--2418
"111110001110010000110001100000000000",--2419
"001111001010000001000000000000000100",--2420
"111110000110001001000001100000000000",--2421
"001011000000000000110000000100101111",--2422
"000101000000000000000000100101111101",--2423
"111110000110100000000001100000000000",--2424
"111110001110000000110001100000000000",--2425
"001111001010000001000000000000000100",--2426
"111110000110001001000001100000000000",--2427
"001011000000000000110000000100101111",--2428
"101001000000000001000000000000000001",--2429
"000101000000000000000000100110000000",--2430
"101000000001111000000010000000000000",--2431
"001111000000000000110000000100101111",--2432
"010000001001000000000000000000101101",--2433
"101111001001110001001011111001001100",--2434
"101111001001100001001100110011001101",--2435
"010110001001000000110000000000101010",--2436
"001101000100000000110000000000000000",--2437
"001001111100000000100000000000000000",--2438
"001001111100000000011111111111111111",--2439
"010011000111000000000000001111110011",--2440
"101111001001110001000011110000100011",--2441
"101111001001100001001101011100001010",--2442
"111110000110000001000001100000000000",--2443
"001111000000000001000000000101100100",--2444
"111110001000001000110010000000000000",--2445
"001111000000000001010000000100101010",--2446
"111110001000000001010010000000000000",--2447
"001111000000000001010000000101100101",--2448
"111110001010001000110010100000000000",--2449
"001111000000000001100000000100101011",--2450
"111110001010000001100010100000000000",--2451
"001111000000000001100000000101100110",--2452
"111110001100001000110001100000000000",--2453
"001111000000000001100000000100101100",--2454
"111110000110000001100001100000000000",--2455
"001101000110000000110000000101101101",--2456
"001101000110000001000000000000000101",--2457
"001111001000000001100000000000000000",--2458
"111110001000010001100011000000000000",--2459
"001111001000000001110000000000000001",--2460
"111110001010010001110011100000000000",--2461
"001111001000000010000000000000000010",--2462
"111110000110010010000100000000000000",--2463
"001101000110000001000000000000000001",--2464
"011111001001000000010000000110000101",--2465
"101110001101111000000011000000000001",--2466
"001101000110000001000000000000000100",--2467
"001111001000000010010000000000000000",--2468
"010110010011000001100000000101111110",--2469
"101110001111111000000011000000000001",--2470
"001111001000000001110000000000000001",--2471
"010110001111000001100000000101111011",--2472
"101110010001111000000011000000000001",--2473
"001111001000000001110000000000000010",--2474
"010110001111000001100000000101111000",--2475
"001101000110000000110000000000000110",--2476
"011100000111000000000000001001011011",--2477
"000101000000000000000000101101011100",--2478
"001101000110000000110000000101101101",--2479
"001101000110000000110000000000000110",--2480
"011100000111000000000000000000000010",--2481
"101000000001111000000000100000000000",--2482
"000100000000000000001111100000000000",--2483
"101001000010000000010000000000000001",--2484
"001100000100000000010001100000000000",--2485
"011111000111000000000000000000000010",--2486
"101000000001111000000000100000000000",--2487
"000100000000000000001111100000000000",--2488
"001100000100000000010001100000000000",--2489
"001101000110000001000000000101101101",--2490
"001111000000000000110000000100101010",--2491
"001101001000000001010000000000000101",--2492
"001111001010000001000000000000000000",--2493
"111110000110010001000001100000000000",--2494
"001111000000000001000000000100101011",--2495
"001111001010000001010000000000000001",--2496
"111110001000010001010010000000000000",--2497
"001111000000000001010000000100101100",--2498
"001111001010000001100000000000000010",--2499
"111110001010010001100010100000000000",--2500
"001101000110000001010000000010111110",--2501
"001101001000000001100000000000000001",--2502
"011111001101000000010000000000111100",--2503
"001111001010000001100000000000000000",--2504
"111110001100010000110011000000000000",--2505
"001111001010000001110000000000000001",--2506
"111110001100001001110011000000000000",--2507
"001111000000000001110000000011111011",--2508
"111110001100001001110011100000000000",--2509
"111110001110000001000011100000000001",--2510
"001101001000000001000000000000000100",--2511
"001111001000000010000000000000000001",--2512
"010110010001000001110000000000000111",--2513
"001111000000000001110000000011111100",--2514
"111110001100001001110011100000000000",--2515
"111110001110000001010011100000000001",--2516
"001111001000000010000000000000000010",--2517
"010110010001000001110000000000000010",--2518
"001111001010000001110000000000000001",--2519
"011110001111000000000000000000101000",--2520
"001111001010000001100000000000000010",--2521
"111110001100010001000011000000000000",--2522
"001111001010000001110000000000000011",--2523
"111110001100001001110011000000000000",--2524
"001111000000000001110000000011111010",--2525
"111110001100001001110011100000000000",--2526
"111110001110000000110011100000000001",--2527
"001111001000000010000000000000000000",--2528
"010110010001000001110000000000000111",--2529
"001111000000000001110000000011111100",--2530
"111110001100001001110011100000000000",--2531
"111110001110000001010011100000000001",--2532
"001111001000000010000000000000000010",--2533
"010110010001000001110000000000000010",--2534
"001111001010000001110000000000000011",--2535
"011110001111000000000000000000010101",--2536
"001111001010000001100000000000000100",--2537
"111110001100010001010010100000000000",--2538
"001111001010000001100000000000000101",--2539
"111110001010001001100010100000000000",--2540
"001111000000000001100000000011111010",--2541
"111110001010001001100011000000000000",--2542
"111110001100000000110001100000000001",--2543
"001111001000000001100000000000000000",--2544
"010110001101000000110000000000000111",--2545
"001111000000000000110000000011111011",--2546
"111110001010001000110001100000000000",--2547
"111110000110000001000001100000000001",--2548
"001111001000000001000000000000000001",--2549
"010110001001000000110000000000000010",--2550
"001111001010000000110000000000000101",--2551
"011110000111000000000000000000000010",--2552
"101000000001111000000010000000000000",--2553
"000101000000000000000000101001010100",--2554
"001011000000000001010000000100101111",--2555
"101001000000000001000000000000000011",--2556
"000101000000000000000000101001010100",--2557
"001011000000000001100000000100101111",--2558
"101001000000000001000000000000000010",--2559
"000101000000000000000000101001010100",--2560
"001011000000000001100000000100101111",--2561
"101001000000000001000000000000000001",--2562
"000101000000000000000000101001010100",--2563
"011111001101000000100000000000001111",--2564
"001111001010000001100000000000000000",--2565
"011010001101000000000000000000001011",--2566
"001111001010000001100000000000000001",--2567
"111110001100001000110001100000000000",--2568
"001111001010000001100000000000000010",--2569
"111110001100001001000010000000000000",--2570
"111110000110000001000001100000000000",--2571
"001111001010000001000000000000000011",--2572
"111110001000001001010010000000000000",--2573
"111110000110000001000001100000000000",--2574
"001011000000000000110000000100101111",--2575
"101001000000000001000000000000000001",--2576
"000101000000000000000000101001010100",--2577
"101000000001111000000010000000000000",--2578
"000101000000000000000000101001010100",--2579
"001111001010000001100000000000000000",--2580
"011110001101000000000000000000000010",--2581
"101000000001111000000010000000000000",--2582
"000101000000000000000000101001010100",--2583
"001111001010000001110000000000000001",--2584
"111110001110001000110011100000000000",--2585
"001111001010000010000000000000000010",--2586
"111110010000001001000100000000000000",--2587
"111110001110000010000011100000000000",--2588
"001111001010000010000000000000000011",--2589
"111110010000001001010100000000000000",--2590
"111110001110000010000011100000000000",--2591
"111110000110001000110100000000000000",--2592
"001101001000000001110000000000000100",--2593
"001111001110000010010000000000000000",--2594
"111110010000001010010100000000000000",--2595
"111110001000001001000100100000000000",--2596
"001111001110000010100000000000000001",--2597
"111110010010001010100100100000000000",--2598
"111110010000000010010100000000000000",--2599
"111110001010001001010100100000000000",--2600
"001111001110000010100000000000000010",--2601
"111110010010001010100100100000000000",--2602
"111110010000000010010100000000000000",--2603
"001101001000000001110000000000000011",--2604
"011100001111000000000000000000000011",--2605
"101110010001111000000001100000000000",--2606
"011111001101000000110000000000010000",--2607
"000101000000000000000000101000111111",--2608
"111110001000001001010100100000000000",--2609
"001101001000000001110000000000001001",--2610
"001111001110000010100000000000000000",--2611
"111110010010001010100100100000000000",--2612
"111110010000000010010100000000000000",--2613
"111110001010001000110010100000000000",--2614
"001111001110000010010000000000000001",--2615
"111110001010001010010010100000000000",--2616
"111110010000000001010010100000000000",--2617
"111110000110001001000001100000000000",--2618
"001111001110000001000000000000000010",--2619
"111110000110001001000001100000000000",--2620
"111110001010000000110001100000000000",--2621
"011111001101000000110000000000000001",--2622
"111110000110010000010001100000000000",--2623
"111110001110001001110010000000000000",--2624
"111110001100001000110001100000000000",--2625
"111110001000010000110001100000000000",--2626
"010110000111000000000000000000001111",--2627
"001101001000000001000000000000000110",--2628
"011100001001000000000000000000000110",--2629
"111110000110100000000001100000000000",--2630
"111110001110010000110001100000000000",--2631
"001111001010000001000000000000000100",--2632
"111110000110001001000001100000000000",--2633
"001011000000000000110000000100101111",--2634
"000101000000000000000000101001010001",--2635
"111110000110100000000001100000000000",--2636
"111110001110000000110001100000000000",--2637
"001111001010000001000000000000000100",--2638
"111110000110001001000001100000000000",--2639
"001011000000000000110000000100101111",--2640
"101001000000000001000000000000000001",--2641
"000101000000000000000000101001010100",--2642
"101000000001111000000010000000000000",--2643
"001111000000000000110000000100101111",--2644
"010000001001000000000000000000101101",--2645
"101111001001110001001011111001001100",--2646
"101111001001100001001100110011001101",--2647
"010110001001000000110000000000101010",--2648
"001101000100000000110000000000000000",--2649
"001001111100000000100000000000000000",--2650
"001001111100000000011111111111111111",--2651
"010011000111000000000000000011000101",--2652
"101111001001110001000011110000100011",--2653
"101111001001100001001101011100001010",--2654
"111110000110000001000001100000000000",--2655
"001111000000000001000000000101100100",--2656
"111110001000001000110010000000000000",--2657
"001111000000000001010000000100101010",--2658
"111110001000000001010010000000000000",--2659
"001111000000000001010000000101100101",--2660
"111110001010001000110010100000000000",--2661
"001111000000000001100000000100101011",--2662
"111110001010000001100010100000000000",--2663
"001111000000000001100000000101100110",--2664
"111110001100001000110001100000000000",--2665
"001111000000000001100000000100101100",--2666
"111110000110000001100001100000000000",--2667
"001101000110000000110000000101101101",--2668
"001101000110000001000000000000000101",--2669
"001111001000000001100000000000000000",--2670
"111110001000010001100011000000000000",--2671
"001111001000000001110000000000000001",--2672
"111110001010010001110011100000000000",--2673
"001111001000000010000000000000000010",--2674
"111110000110010010000100000000000000",--2675
"001101000110000001000000000000000001",--2676
"011111001001000000010000000000010111",--2677
"101110001101111000000011000000000001",--2678
"001101000110000001000000000000000100",--2679
"001111001000000010010000000000000000",--2680
"010110010011000001100000000000010000",--2681
"101110001111111000000011000000000001",--2682
"001111001000000001110000000000000001",--2683
"010110001111000001100000000000001101",--2684
"101110010001111000000011000000000001",--2685
"001111001000000001110000000000000010",--2686
"010110001111000001100000000000001010",--2687
"001101000110000000110000000000000110",--2688
"011100000111000000000000000010011100",--2689
"000101000000000000000000101011000010",--2690
"001101000110000000110000000101101101",--2691
"001101000110000000110000000000000110",--2692
"011100000111000000000000000000000010",--2693
"101000000001111000000000100000000000",--2694
"000100000000000000001111100000000000",--2695
"101001000010000000010000000000000001",--2696
"000101000000000000000000100011100001",--2697
"001101000110000000110000000000000110",--2698
"011100000111000000000000000000110110",--2699
"000101000000000000000000101100011110",--2700
"011111001001000000100000000000001111",--2701
"001101000110000001000000000000000100",--2702
"001111001000000010010000000000000000",--2703
"111110010010001001100011000000000000",--2704
"001111001000000010010000000000000001",--2705
"111110010010001001110011100000000000",--2706
"111110001100000001110011000000000000",--2707
"001111001000000001110000000000000010",--2708
"111110001110001010000011100000000000",--2709
"111110001100000001110011000000000000",--2710
"001101000110000000110000000000000110",--2711
"011010001101000000000000000000000010",--2712
"011111000111000000010000000000101000",--2713
"000101000000000000000000101100011110",--2714
"011100000111000000000000000000100110",--2715
"000101000000000000000000101100011110",--2716
"111110001100001001100100100000000000",--2717
"001101000110000001010000000000000100",--2718
"001111001010000010100000000000000000",--2719
"111110010010001010100100100000000000",--2720
"111110001110001001110101000000000000",--2721
"001111001010000010110000000000000001",--2722
"111110010100001010110101000000000000",--2723
"111110010010000010100100100000000000",--2724
"111110010000001010000101000000000000",--2725
"001111001010000010110000000000000010",--2726
"111110010100001010110101000000000000",--2727
"111110010010000010100100100000000000",--2728
"001101000110000001010000000000000011",--2729
"011100001011000000000000000000000011",--2730
"101110010011111000000011000000000000",--2731
"011111001001000000110000000000010000",--2732
"000101000000000000000000101010111100",--2733
"111110001110001010000101000000000000",--2734
"001101000110000001010000000000001001",--2735
"001111001010000010110000000000000000",--2736
"111110010100001010110101000000000000",--2737
"111110010010000010100100100000000000",--2738
"111110010000001001100100000000000000",--2739
"001111001010000010100000000000000001",--2740
"111110010000001010100100000000000000",--2741
"111110010010000010000100000000000000",--2742
"111110001100001001110011000000000000",--2743
"001111001010000001110000000000000010",--2744
"111110001100001001110011000000000000",--2745
"111110010000000001100011000000000000",--2746
"011111001001000000110000000000000001",--2747
"111110001100010000010011000000000000",--2748
"001101000110000000110000000000000110",--2749
"011010001101000000000000000000000010",--2750
"011111000111000000010000000000000010",--2751
"000101000000000000000000101100011110",--2752
"010000000111000000000000000001011100",--2753
"001101000100000000110000000000000001",--2754
"010011000111000000000000000001011110",--2755
"001101000110000000110000000101101101",--2756
"001101000110000001000000000000000101",--2757
"001111001000000001100000000000000000",--2758
"111110001000010001100011000000000000",--2759
"001111001000000001110000000000000001",--2760
"111110001010010001110011100000000000",--2761
"001111001000000010000000000000000010",--2762
"111110000110010010000100000000000000",--2763
"001101000110000001000000000000000001",--2764
"011111001001000000010000000000010000",--2765
"101110001101111000000011000000000001",--2766
"001101000110000001000000000000000100",--2767
"001111001000000010010000000000000000",--2768
"010110010011000001100000000000001001",--2769
"101110001111111000000011000000000001",--2770
"001111001000000001110000000000000001",--2771
"010110001111000001100000000000000110",--2772
"101110010001111000000011000000000001",--2773
"001111001000000001110000000000000010",--2774
"010110001111000001100000000000000011",--2775
"001101000110000000110000000000000110",--2776
"011100000111000000000000000001000100",--2777
"000101000000000000000000101100010011",--2778
"001101000110000000110000000000000110",--2779
"011100000111000000000000000000110110",--2780
"000101000000000000000000101100011110",--2781
"011111001001000000100000000000001111",--2782
"001101000110000001000000000000000100",--2783
"001111001000000010010000000000000000",--2784
"111110010010001001100011000000000000",--2785
"001111001000000010010000000000000001",--2786
"111110010010001001110011100000000000",--2787
"111110001100000001110011000000000000",--2788
"001111001000000001110000000000000010",--2789
"111110001110001010000011100000000000",--2790
"111110001100000001110011000000000000",--2791
"001101000110000000110000000000000110",--2792
"011010001101000000000000000000000010",--2793
"011111000111000000010000000000101000",--2794
"000101000000000000000000101100011110",--2795
"011100000111000000000000000000100110",--2796
"000101000000000000000000101100011110",--2797
"111110001100001001100100100000000000",--2798
"001101000110000001010000000000000100",--2799
"001111001010000010100000000000000000",--2800
"111110010010001010100100100000000000",--2801
"111110001110001001110101000000000000",--2802
"001111001010000010110000000000000001",--2803
"111110010100001010110101000000000000",--2804
"111110010010000010100100100000000000",--2805
"111110010000001010000101000000000000",--2806
"001111001010000010110000000000000010",--2807
"111110010100001010110101000000000000",--2808
"111110010010000010100100100000000000",--2809
"001101000110000001010000000000000011",--2810
"011100001011000000000000000000000011",--2811
"101110010011111000000011000000000000",--2812
"011111001001000000110000000000010000",--2813
"000101000000000000000000101100001101",--2814
"111110001110001010000101000000000000",--2815
"001101000110000001010000000000001001",--2816
"001111001010000010110000000000000000",--2817
"111110010100001010110101000000000000",--2818
"111110010010000010100100100000000000",--2819
"111110010000001001100100000000000000",--2820
"001111001010000010100000000000000001",--2821
"111110010000001010100100000000000000",--2822
"111110010010000010000100000000000000",--2823
"111110001100001001110011000000000000",--2824
"001111001010000001110000000000000010",--2825
"111110001100001001110011000000000000",--2826
"111110010000000001100011000000000000",--2827
"011111001001000000110000000000000001",--2828
"111110001100010000010011000000000000",--2829
"001101000110000000110000000000000110",--2830
"011010001101000000000000000000000010",--2831
"011111000111000000010000000000000010",--2832
"000101000000000000000000101100011110",--2833
"010000000111000000000000000000001011",--2834
"101001000000000000010000000000000010",--2835
"101110001011111000001111100000000000",--2836
"101110000111111000000010100000000000",--2837
"101110001001111000000001100000000000",--2838
"101110111111111000000010000000000000",--2839
"001001111100000111111111111111111110",--2840
"101001111100010111100000000000000011",--2841
"000111000000000000000000011110001000",--2842
"101001111100000111100000000000000011",--2843
"001101111100000111111111111111111110",--2844
"011100000011000000000000000000000100",--2845
"001101111100000000011111111111111111",--2846
"101001000010000000010000000000000001",--2847
"001101111100000000100000000000000000",--2848
"000101000000000000000000100011100001",--2849
"101001000000000000010000000000000001",--2850
"000100000000000000001111100000000000",--2851
"001101000110000000110000000000000110",--2852
"011100000111000000000000000000110110",--2853
"000101000000000000000000110000001001",--2854
"011111001001000000100000000000001111",--2855
"001101000110000001000000000000000100",--2856
"001111001000000010010000000000000000",--2857
"111110010010001001100011000000000000",--2858
"001111001000000010010000000000000001",--2859
"111110010010001001110011100000000000",--2860
"111110001100000001110011000000000000",--2861
"001111001000000001110000000000000010",--2862
"111110001110001010000011100000000000",--2863
"111110001100000001110011000000000000",--2864
"001101000110000000110000000000000110",--2865
"011010001101000000000000000000000010",--2866
"011111000111000000010000000000101000",--2867
"000101000000000000000000110000001001",--2868
"011100000111000000000000000000100110",--2869
"000101000000000000000000110000001001",--2870
"111110001100001001100100100000000000",--2871
"001101000110000001010000000000000100",--2872
"001111001010000010100000000000000000",--2873
"111110010010001010100100100000000000",--2874
"111110001110001001110101000000000000",--2875
"001111001010000010110000000000000001",--2876
"111110010100001010110101000000000000",--2877
"111110010010000010100100100000000000",--2878
"111110010000001010000101000000000000",--2879
"001111001010000010110000000000000010",--2880
"111110010100001010110101000000000000",--2881
"111110010010000010100100100000000000",--2882
"001101000110000001010000000000000011",--2883
"011100001011000000000000000000000011",--2884
"101110010011111000000011000000000000",--2885
"011111001001000000110000000000010000",--2886
"000101000000000000000000101101010110",--2887
"111110001110001010000101000000000000",--2888
"001101000110000001010000000000001001",--2889
"001111001010000010110000000000000000",--2890
"111110010100001010110101000000000000",--2891
"111110010010000010100100100000000000",--2892
"111110010000001001100100000000000000",--2893
"001111001010000010100000000000000001",--2894
"111110010000001010100100000000000000",--2895
"111110010010000010000100000000000000",--2896
"111110001100001001110011000000000000",--2897
"001111001010000001110000000000000010",--2898
"111110001100001001110011000000000000",--2899
"111110010000000001100011000000000000",--2900
"011111001001000000110000000000000001",--2901
"111110001100010000010011000000000000",--2902
"001101000110000000110000000000000110",--2903
"011010001101000000000000000000000010",--2904
"011111000111000000010000000000000010",--2905
"000101000000000000000000110000001001",--2906
"010000000111000000000000000010101101",--2907
"001101000100000000110000000000000001",--2908
"010011000111000000000000001000011110",--2909
"001101000110000000110000000101101101",--2910
"001101000110000001000000000000000101",--2911
"001111001000000001100000000000000000",--2912
"111110001000010001100011000000000000",--2913
"001111001000000001110000000000000001",--2914
"111110001010010001110011100000000000",--2915
"001111001000000010000000000000000010",--2916
"111110000110010010000100000000000000",--2917
"001101000110000001000000000000000001",--2918
"011111001001000000010000000000010000",--2919
"101110001101111000000011000000000001",--2920
"001101000110000001000000000000000100",--2921
"001111001000000010010000000000000000",--2922
"010110010011000001100000000000001001",--2923
"101110001111111000000011000000000001",--2924
"001111001000000001110000000000000001",--2925
"010110001111000001100000000000000110",--2926
"101110010001111000000011000000000001",--2927
"001111001000000001110000000000000010",--2928
"010110001111000001100000000000000011",--2929
"001101000110000000110000000000000110",--2930
"011100000111000000000000000010010101",--2931
"000101000000000000000000101110101101",--2932
"001101000110000000110000000000000110",--2933
"011100000111000000000000000000110110",--2934
"000101000000000000000000110000001001",--2935
"011111001001000000100000000000001111",--2936
"001101000110000001000000000000000100",--2937
"001111001000000010010000000000000000",--2938
"111110010010001001100011000000000000",--2939
"001111001000000010010000000000000001",--2940
"111110010010001001110011100000000000",--2941
"111110001100000001110011000000000000",--2942
"001111001000000001110000000000000010",--2943
"111110001110001010000011100000000000",--2944
"111110001100000001110011000000000000",--2945
"001101000110000000110000000000000110",--2946
"011010001101000000000000000000000010",--2947
"011111000111000000010000000000101000",--2948
"000101000000000000000000110000001001",--2949
"011100000111000000000000000000100110",--2950
"000101000000000000000000110000001001",--2951
"111110001100001001100100100000000000",--2952
"001101000110000001010000000000000100",--2953
"001111001010000010100000000000000000",--2954
"111110010010001010100100100000000000",--2955
"111110001110001001110101000000000000",--2956
"001111001010000010110000000000000001",--2957
"111110010100001010110101000000000000",--2958
"111110010010000010100100100000000000",--2959
"111110010000001010000101000000000000",--2960
"001111001010000010110000000000000010",--2961
"111110010100001010110101000000000000",--2962
"111110010010000010100100100000000000",--2963
"001101000110000001010000000000000011",--2964
"011100001011000000000000000000000011",--2965
"101110010011111000000011000000000000",--2966
"011111001001000000110000000000010000",--2967
"000101000000000000000000101110100111",--2968
"111110001110001010000101000000000000",--2969
"001101000110000001010000000000001001",--2970
"001111001010000010110000000000000000",--2971
"111110010100001010110101000000000000",--2972
"111110010010000010100100100000000000",--2973
"111110010000001001100100000000000000",--2974
"001111001010000010100000000000000001",--2975
"111110010000001010100100000000000000",--2976
"111110010010000010000100000000000000",--2977
"111110001100001001110011000000000000",--2978
"001111001010000001110000000000000010",--2979
"111110001100001001110011000000000000",--2980
"111110010000000001100011000000000000",--2981
"011111001001000000110000000000000001",--2982
"111110001100010000010011000000000000",--2983
"001101000110000000110000000000000110",--2984
"011010001101000000000000000000000010",--2985
"011111000111000000010000000000000010",--2986
"000101000000000000000000110000001001",--2987
"010000000111000000000000000001011100",--2988
"001101000100000000110000000000000010",--2989
"010011000111000000000000000111001101",--2990
"001101000110000000110000000101101101",--2991
"001101000110000001000000000000000101",--2992
"001111001000000001100000000000000000",--2993
"111110001000010001100011000000000000",--2994
"001111001000000001110000000000000001",--2995
"111110001010010001110011100000000000",--2996
"001111001000000010000000000000000010",--2997
"111110000110010010000100000000000000",--2998
"001101000110000001000000000000000001",--2999
"011111001001000000010000000000010000",--3000
"101110001101111000000011000000000001",--3001
"001101000110000001000000000000000100",--3002
"001111001000000010010000000000000000",--3003
"010110010011000001100000000000001001",--3004
"101110001111111000000011000000000001",--3005
"001111001000000001110000000000000001",--3006
"010110001111000001100000000000000110",--3007
"101110010001111000000011000000000001",--3008
"001111001000000001110000000000000010",--3009
"010110001111000001100000000000000011",--3010
"001101000110000000110000000000000110",--3011
"011100000111000000000000000001000100",--3012
"000101000000000000000000101111111110",--3013
"001101000110000000110000000000000110",--3014
"011100000111000000000000000000110110",--3015
"000101000000000000000000110000001001",--3016
"011111001001000000100000000000001111",--3017
"001101000110000001000000000000000100",--3018
"001111001000000010010000000000000000",--3019
"111110010010001001100011000000000000",--3020
"001111001000000010010000000000000001",--3021
"111110010010001001110011100000000000",--3022
"111110001100000001110011000000000000",--3023
"001111001000000001110000000000000010",--3024
"111110001110001010000011100000000000",--3025
"111110001100000001110011000000000000",--3026
"001101000110000000110000000000000110",--3027
"011010001101000000000000000000000010",--3028
"011111000111000000010000000000101000",--3029
"000101000000000000000000110000001001",--3030
"011100000111000000000000000000100110",--3031
"000101000000000000000000110000001001",--3032
"111110001100001001100100100000000000",--3033
"001101000110000001010000000000000100",--3034
"001111001010000010100000000000000000",--3035
"111110010010001010100100100000000000",--3036
"111110001110001001110101000000000000",--3037
"001111001010000010110000000000000001",--3038
"111110010100001010110101000000000000",--3039
"111110010010000010100100100000000000",--3040
"111110010000001010000101000000000000",--3041
"001111001010000010110000000000000010",--3042
"111110010100001010110101000000000000",--3043
"111110010010000010100100100000000000",--3044
"001101000110000001010000000000000011",--3045
"011100001011000000000000000000000011",--3046
"101110010011111000000011000000000000",--3047
"011111001001000000110000000000010000",--3048
"000101000000000000000000101111111000",--3049
"111110001110001010000101000000000000",--3050
"001101000110000001010000000000001001",--3051
"001111001010000010110000000000000000",--3052
"111110010100001010110101000000000000",--3053
"111110010010000010100100100000000000",--3054
"111110010000001001100100000000000000",--3055
"001111001010000010100000000000000001",--3056
"111110010000001010100100000000000000",--3057
"111110010010000010000100000000000000",--3058
"111110001100001001110011000000000000",--3059
"001111001010000001110000000000000010",--3060
"111110001100001001110011000000000000",--3061
"111110010000000001100011000000000000",--3062
"011111001001000000110000000000000001",--3063
"111110001100010000010011000000000000",--3064
"001101000110000000110000000000000110",--3065
"011010001101000000000000000000000010",--3066
"011111000111000000010000000000000010",--3067
"000101000000000000000000110000001001",--3068
"010000000111000000000000000000001011",--3069
"101001000000000000010000000000000011",--3070
"101110001011111000001111100000000000",--3071
"101110000111111000000010100000000000",--3072
"101110001001111000000001100000000000",--3073
"101110111111111000000010000000000000",--3074
"001001111100000111111111111111111110",--3075
"101001111100010111100000000000000011",--3076
"000111000000000000000000011110001000",--3077
"101001111100000111100000000000000011",--3078
"001101111100000111111111111111111110",--3079
"011100000011000000000000000101110011",--3080
"001101111100000000011111111111111111",--3081
"101001000010000000010000000000000001",--3082
"001101111100000000110000000000000000",--3083
"001100000110000000010001000000000000",--3084
"011111000101000000000000000000000010",--3085
"101000000001111000000000100000000000",--3086
"000100000000000000001111100000000000",--3087
"001100000110000000010001000000000000",--3088
"001101000100000001000000000101101101",--3089
"001111000000000000110000000100101010",--3090
"001101001000000001010000000000000101",--3091
"001111001010000001000000000000000000",--3092
"111110000110010001000001100000000000",--3093
"001111000000000001000000000100101011",--3094
"001111001010000001010000000000000001",--3095
"111110001000010001010010000000000000",--3096
"001111000000000001010000000100101100",--3097
"001111001010000001100000000000000010",--3098
"111110001010010001100010100000000000",--3099
"001101000100000001010000000010111110",--3100
"001101001000000001100000000000000001",--3101
"011111001101000000010000000000111100",--3102
"001111001010000001100000000000000000",--3103
"111110001100010000110011000000000000",--3104
"001111001010000001110000000000000001",--3105
"111110001100001001110011000000000000",--3106
"001111000000000001110000000011111011",--3107
"111110001100001001110011100000000000",--3108
"111110001110000001000011100000000001",--3109
"001101001000000001000000000000000100",--3110
"001111001000000010000000000000000001",--3111
"010110010001000001110000000000000111",--3112
"001111000000000001110000000011111100",--3113
"111110001100001001110011100000000000",--3114
"111110001110000001010011100000000001",--3115
"001111001000000010000000000000000010",--3116
"010110010001000001110000000000000010",--3117
"001111001010000001110000000000000001",--3118
"011110001111000000000000000000101000",--3119
"001111001010000001100000000000000010",--3120
"111110001100010001000011000000000000",--3121
"001111001010000001110000000000000011",--3122
"111110001100001001110011000000000000",--3123
"001111000000000001110000000011111010",--3124
"111110001100001001110011100000000000",--3125
"111110001110000000110011100000000001",--3126
"001111001000000010000000000000000000",--3127
"010110010001000001110000000000000111",--3128
"001111000000000001110000000011111100",--3129
"111110001100001001110011100000000000",--3130
"111110001110000001010011100000000001",--3131
"001111001000000010000000000000000010",--3132
"010110010001000001110000000000000010",--3133
"001111001010000001110000000000000011",--3134
"011110001111000000000000000000010101",--3135
"001111001010000001100000000000000100",--3136
"111110001100010001010010100000000000",--3137
"001111001010000001100000000000000101",--3138
"111110001010001001100010100000000000",--3139
"001111000000000001100000000011111010",--3140
"111110001010001001100011000000000000",--3141
"111110001100000000110001100000000001",--3142
"001111001000000001100000000000000000",--3143
"010110001101000000110000000000000111",--3144
"001111000000000000110000000011111011",--3145
"111110001010001000110001100000000000",--3146
"111110000110000001000001100000000001",--3147
"001111001000000001000000000000000001",--3148
"010110001001000000110000000000000010",--3149
"001111001010000000110000000000000101",--3150
"011110000111000000000000000000000010",--3151
"101000000001111000000010000000000000",--3152
"000101000000000000000000110010101011",--3153
"001011000000000001010000000100101111",--3154
"101001000000000001000000000000000011",--3155
"000101000000000000000000110010101011",--3156
"001011000000000001100000000100101111",--3157
"101001000000000001000000000000000010",--3158
"000101000000000000000000110010101011",--3159
"001011000000000001100000000100101111",--3160
"101001000000000001000000000000000001",--3161
"000101000000000000000000110010101011",--3162
"011111001101000000100000000000001111",--3163
"001111001010000001100000000000000000",--3164
"011010001101000000000000000000001011",--3165
"001111001010000001100000000000000001",--3166
"111110001100001000110001100000000000",--3167
"001111001010000001100000000000000010",--3168
"111110001100001001000010000000000000",--3169
"111110000110000001000001100000000000",--3170
"001111001010000001000000000000000011",--3171
"111110001000001001010010000000000000",--3172
"111110000110000001000001100000000000",--3173
"001011000000000000110000000100101111",--3174
"101001000000000001000000000000000001",--3175
"000101000000000000000000110010101011",--3176
"101000000001111000000010000000000000",--3177
"000101000000000000000000110010101011",--3178
"001111001010000001100000000000000000",--3179
"011110001101000000000000000000000010",--3180
"101000000001111000000010000000000000",--3181
"000101000000000000000000110010101011",--3182
"001111001010000001110000000000000001",--3183
"111110001110001000110011100000000000",--3184
"001111001010000010000000000000000010",--3185
"111110010000001001000100000000000000",--3186
"111110001110000010000011100000000000",--3187
"001111001010000010000000000000000011",--3188
"111110010000001001010100000000000000",--3189
"111110001110000010000011100000000000",--3190
"111110000110001000110100000000000000",--3191
"001101001000000001110000000000000100",--3192
"001111001110000010010000000000000000",--3193
"111110010000001010010100000000000000",--3194
"111110001000001001000100100000000000",--3195
"001111001110000010100000000000000001",--3196
"111110010010001010100100100000000000",--3197
"111110010000000010010100000000000000",--3198
"111110001010001001010100100000000000",--3199
"001111001110000010100000000000000010",--3200
"111110010010001010100100100000000000",--3201
"111110010000000010010100000000000000",--3202
"001101001000000001110000000000000011",--3203
"011100001111000000000000000000000011",--3204
"101110010001111000000001100000000000",--3205
"011111001101000000110000000000010000",--3206
"000101000000000000000000110010010110",--3207
"111110001000001001010100100000000000",--3208
"001101001000000001110000000000001001",--3209
"001111001110000010100000000000000000",--3210
"111110010010001010100100100000000000",--3211
"111110010000000010010100000000000000",--3212
"111110001010001000110010100000000000",--3213
"001111001110000010010000000000000001",--3214
"111110001010001010010010100000000000",--3215
"111110010000000001010010100000000000",--3216
"111110000110001001000001100000000000",--3217
"001111001110000001000000000000000010",--3218
"111110000110001001000001100000000000",--3219
"111110001010000000110001100000000000",--3220
"011111001101000000110000000000000001",--3221
"111110000110010000010001100000000000",--3222
"111110001110001001110010000000000000",--3223
"111110001100001000110001100000000000",--3224
"111110001000010000110001100000000000",--3225
"010110000111000000000000000000001111",--3226
"001101001000000001000000000000000110",--3227
"011100001001000000000000000000000110",--3228
"111110000110100000000001100000000000",--3229
"111110001110010000110001100000000000",--3230
"001111001010000001000000000000000100",--3231
"111110000110001001000001100000000000",--3232
"001011000000000000110000000100101111",--3233
"000101000000000000000000110010101000",--3234
"111110000110100000000001100000000000",--3235
"111110001110000000110001100000000000",--3236
"001111001010000001000000000000000100",--3237
"111110000110001001000001100000000000",--3238
"001011000000000000110000000100101111",--3239
"101001000000000001000000000000000001",--3240
"000101000000000000000000110010101011",--3241
"101000000001111000000010000000000000",--3242
"001111000000000000110000000100101111",--3243
"010000001001000000000000000000101100",--3244
"101111001001110001001011111001001100",--3245
"101111001001100001001100110011001101",--3246
"010110001001000000110000000000101001",--3247
"001101000110000000100000000000000000",--3248
"001001111100000000011111111111111110",--3249
"010011000101000000000000000011000111",--3250
"101111001001110001000011110000100011",--3251
"101111001001100001001101011100001010",--3252
"111110000110000001000001100000000000",--3253
"001111000000000001000000000101100100",--3254
"111110001000001000110010000000000000",--3255
"001111000000000001010000000100101010",--3256
"111110001000000001010010000000000000",--3257
"001111000000000001010000000101100101",--3258
"111110001010001000110010100000000000",--3259
"001111000000000001100000000100101011",--3260
"111110001010000001100010100000000000",--3261
"001111000000000001100000000101100110",--3262
"111110001100001000110001100000000000",--3263
"001111000000000001100000000100101100",--3264
"111110000110000001100001100000000000",--3265
"001101000100000000100000000101101101",--3266
"001101000100000001000000000000000101",--3267
"001111001000000001100000000000000000",--3268
"111110001000010001100011000000000000",--3269
"001111001000000001110000000000000001",--3270
"111110001010010001110011100000000000",--3271
"001111001000000010000000000000000010",--3272
"111110000110010010000100000000000000",--3273
"001101000100000001000000000000000001",--3274
"011111001001000000010000000000011000",--3275
"101110001101111000000011000000000001",--3276
"001101000100000001000000000000000100",--3277
"001111001000000010010000000000000000",--3278
"010110010011000001100000000000010001",--3279
"101110001111111000000011000000000001",--3280
"001111001000000001110000000000000001",--3281
"010110001111000001100000000000001110",--3282
"101110010001111000000011000000000001",--3283
"001111001000000001110000000000000010",--3284
"010110001111000001100000000000001011",--3285
"001101000100000000100000000000000110",--3286
"011100000101000000000000000010011110",--3287
"000101000000000000000000110100011001",--3288
"001101000100000000100000000101101101",--3289
"001101000100000000100000000000000110",--3290
"011100000101000000000000000000000010",--3291
"101000000001111000000000100000000000",--3292
"000100000000000000001111100000000000",--3293
"101001000010000000010000000000000001",--3294
"101000000111111000000001000000000000",--3295
"000101000000000000000000100011100001",--3296
"001101000100000000100000000000000110",--3297
"011100000101000000000000000000110110",--3298
"000101000000000000000000110101110110",--3299
"011111001001000000100000000000001111",--3300
"001101000100000001000000000000000100",--3301
"001111001000000010010000000000000000",--3302
"111110010010001001100011000000000000",--3303
"001111001000000010010000000000000001",--3304
"111110010010001001110011100000000000",--3305
"111110001100000001110011000000000000",--3306
"001111001000000001110000000000000010",--3307
"111110001110001010000011100000000000",--3308
"111110001100000001110011000000000000",--3309
"001101000100000000100000000000000110",--3310
"011010001101000000000000000000000010",--3311
"011111000101000000010000000000101000",--3312
"000101000000000000000000110101110110",--3313
"011100000101000000000000000000100110",--3314
"000101000000000000000000110101110110",--3315
"111110001100001001100100100000000000",--3316
"001101000100000001010000000000000100",--3317
"001111001010000010100000000000000000",--3318
"111110010010001010100100100000000000",--3319
"111110001110001001110101000000000000",--3320
"001111001010000010110000000000000001",--3321
"111110010100001010110101000000000000",--3322
"111110010010000010100100100000000000",--3323
"111110010000001010000101000000000000",--3324
"001111001010000010110000000000000010",--3325
"111110010100001010110101000000000000",--3326
"111110010010000010100100100000000000",--3327
"001101000100000001010000000000000011",--3328
"011100001011000000000000000000000011",--3329
"101110010011111000000011000000000000",--3330
"011111001001000000110000000000010000",--3331
"000101000000000000000000110100010011",--3332
"111110001110001010000101000000000000",--3333
"001101000100000001010000000000001001",--3334
"001111001010000010110000000000000000",--3335
"111110010100001010110101000000000000",--3336
"111110010010000010100100100000000000",--3337
"111110010000001001100100000000000000",--3338
"001111001010000010100000000000000001",--3339
"111110010000001010100100000000000000",--3340
"111110010010000010000100000000000000",--3341
"111110001100001001110011000000000000",--3342
"001111001010000001110000000000000010",--3343
"111110001100001001110011000000000000",--3344
"111110010000000001100011000000000000",--3345
"011111001001000000110000000000000001",--3346
"111110001100010000010011000000000000",--3347
"001101000100000000100000000000000110",--3348
"011010001101000000000000000000000010",--3349
"011111000101000000010000000000000010",--3350
"000101000000000000000000110101110110",--3351
"010000000101000000000000000001011101",--3352
"001101000110000000100000000000000001",--3353
"010011000101000000000000000001011111",--3354
"001101000100000000100000000101101101",--3355
"001101000100000001000000000000000101",--3356
"001111001000000001100000000000000000",--3357
"111110001000010001100011000000000000",--3358
"001111001000000001110000000000000001",--3359
"111110001010010001110011100000000000",--3360
"001111001000000010000000000000000010",--3361
"111110000110010010000100000000000000",--3362
"001101000100000001000000000000000001",--3363
"011111001001000000010000000000010000",--3364
"101110001101111000000011000000000001",--3365
"001101000100000001000000000000000100",--3366
"001111001000000010010000000000000000",--3367
"010110010011000001100000000000001001",--3368
"101110001111111000000011000000000001",--3369
"001111001000000001110000000000000001",--3370
"010110001111000001100000000000000110",--3371
"101110010001111000000011000000000001",--3372
"001111001000000001110000000000000010",--3373
"010110001111000001100000000000000011",--3374
"001101000100000000100000000000000110",--3375
"011100000101000000000000000001000101",--3376
"000101000000000000000000110101101010",--3377
"001101000100000000100000000000000110",--3378
"011100000101000000000000000000110110",--3379
"000101000000000000000000110101110110",--3380
"011111001001000000100000000000001111",--3381
"001101000100000001000000000000000100",--3382
"001111001000000010010000000000000000",--3383
"111110010010001001100011000000000000",--3384
"001111001000000010010000000000000001",--3385
"111110010010001001110011100000000000",--3386
"111110001100000001110011000000000000",--3387
"001111001000000001110000000000000010",--3388
"111110001110001010000011100000000000",--3389
"111110001100000001110011000000000000",--3390
"001101000100000000100000000000000110",--3391
"011010001101000000000000000000000010",--3392
"011111000101000000010000000000101000",--3393
"000101000000000000000000110101110110",--3394
"011100000101000000000000000000100110",--3395
"000101000000000000000000110101110110",--3396
"111110001100001001100100100000000000",--3397
"001101000100000001010000000000000100",--3398
"001111001010000010100000000000000000",--3399
"111110010010001010100100100000000000",--3400
"111110001110001001110101000000000000",--3401
"001111001010000010110000000000000001",--3402
"111110010100001010110101000000000000",--3403
"111110010010000010100100100000000000",--3404
"111110010000001010000101000000000000",--3405
"001111001010000010110000000000000010",--3406
"111110010100001010110101000000000000",--3407
"111110010010000010100100100000000000",--3408
"001101000100000001010000000000000011",--3409
"011100001011000000000000000000000011",--3410
"101110010011111000000011000000000000",--3411
"011111001001000000110000000000010000",--3412
"000101000000000000000000110101100100",--3413
"111110001110001010000101000000000000",--3414
"001101000100000001010000000000001001",--3415
"001111001010000010110000000000000000",--3416
"111110010100001010110101000000000000",--3417
"111110010010000010100100100000000000",--3418
"111110010000001001100100000000000000",--3419
"001111001010000010100000000000000001",--3420
"111110010000001010100100000000000000",--3421
"111110010010000010000100000000000000",--3422
"111110001100001001110011000000000000",--3423
"001111001010000001110000000000000010",--3424
"111110001100001001110011000000000000",--3425
"111110010000000001100011000000000000",--3426
"011111001001000000110000000000000001",--3427
"111110001100010000010011000000000000",--3428
"001101000100000000100000000000000110",--3429
"011010001101000000000000000000000010",--3430
"011111000101000000010000000000000010",--3431
"000101000000000000000000110101110110",--3432
"010000000101000000000000000000001100",--3433
"101001000000000000010000000000000010",--3434
"101000000111111000000001000000000000",--3435
"101110001011111000001111100000000000",--3436
"101110000111111000000010100000000000",--3437
"101110001001111000000001100000000000",--3438
"101110111111111000000010000000000000",--3439
"001001111100000111111111111111111101",--3440
"101001111100010111100000000000000100",--3441
"000111000000000000000000011110001000",--3442
"101001111100000111100000000000000100",--3443
"001101111100000111111111111111111101",--3444
"011100000011000000000000000000000100",--3445
"001101111100000000011111111111111110",--3446
"101001000010000000010000000000000001",--3447
"001101111100000000100000000000000000",--3448
"000101000000000000000000100011100001",--3449
"101001000000000000010000000000000001",--3450
"000100000000000000001111100000000000",--3451
"101001000000000000010000000000000001",--3452
"000100000000000000001111100000000000",--3453
"001100000100000000010001100000000000",--3454
"011111000111000000000000000000000010",--3455
"101000000001111000000000100000000000",--3456
"000100000000000000001111100000000000",--3457
"001101000110000000110000000100110001",--3458
"001101000110000001000000000000000000",--3459
"001001111100000000100000000000000000",--3460
"001001111100000000011111111111111111",--3461
"010011001001000000000000000101110001",--3462
"001101001000000001010000000101101101",--3463
"001111000000000000110000000100101010",--3464
"001101001010000001100000000000000101",--3465
"001111001100000001000000000000000000",--3466
"111110000110010001000001100000000000",--3467
"001111000000000001000000000100101011",--3468
"001111001100000001010000000000000001",--3469
"111110001000010001010010000000000000",--3470
"001111000000000001010000000100101100",--3471
"001111001100000001100000000000000010",--3472
"111110001010010001100010100000000000",--3473
"001101001000000001100000000010111110",--3474
"001101001010000001110000000000000001",--3475
"011111001111000000010000000000111100",--3476
"001111001100000001100000000000000000",--3477
"111110001100010000110011000000000000",--3478
"001111001100000001110000000000000001",--3479
"111110001100001001110011000000000000",--3480
"001111000000000001110000000011111011",--3481
"111110001100001001110011100000000000",--3482
"111110001110000001000011100000000001",--3483
"001101001010000001010000000000000100",--3484
"001111001010000010000000000000000001",--3485
"010110010001000001110000000000000111",--3486
"001111000000000001110000000011111100",--3487
"111110001100001001110011100000000000",--3488
"111110001110000001010011100000000001",--3489
"001111001010000010000000000000000010",--3490
"010110010001000001110000000000000010",--3491
"001111001100000001110000000000000001",--3492
"011110001111000000000000000000101000",--3493
"001111001100000001100000000000000010",--3494
"111110001100010001000011000000000000",--3495
"001111001100000001110000000000000011",--3496
"111110001100001001110011000000000000",--3497
"001111000000000001110000000011111010",--3498
"111110001100001001110011100000000000",--3499
"111110001110000000110011100000000001",--3500
"001111001010000010000000000000000000",--3501
"010110010001000001110000000000000111",--3502
"001111000000000001110000000011111100",--3503
"111110001100001001110011100000000000",--3504
"111110001110000001010011100000000001",--3505
"001111001010000010000000000000000010",--3506
"010110010001000001110000000000000010",--3507
"001111001100000001110000000000000011",--3508
"011110001111000000000000000000010101",--3509
"001111001100000001100000000000000100",--3510
"111110001100010001010010100000000000",--3511
"001111001100000001100000000000000101",--3512
"111110001010001001100010100000000000",--3513
"001111000000000001100000000011111010",--3514
"111110001010001001100011000000000000",--3515
"111110001100000000110001100000000001",--3516
"001111001010000001100000000000000000",--3517
"010110001101000000110000000000000111",--3518
"001111000000000000110000000011111011",--3519
"111110001010001000110001100000000000",--3520
"111110000110000001000001100000000001",--3521
"001111001010000001000000000000000001",--3522
"010110001001000000110000000000000010",--3523
"001111001100000000110000000000000101",--3524
"011110000111000000000000000000000010",--3525
"101000000001111000000010100000000000",--3526
"000101000000000000000000111000100001",--3527
"001011000000000001010000000100101111",--3528
"101001000000000001010000000000000011",--3529
"000101000000000000000000111000100001",--3530
"001011000000000001100000000100101111",--3531
"101001000000000001010000000000000010",--3532
"000101000000000000000000111000100001",--3533
"001011000000000001100000000100101111",--3534
"101001000000000001010000000000000001",--3535
"000101000000000000000000111000100001",--3536
"011111001111000000100000000000001111",--3537
"001111001100000001100000000000000000",--3538
"011010001101000000000000000000001011",--3539
"001111001100000001100000000000000001",--3540
"111110001100001000110001100000000000",--3541
"001111001100000001100000000000000010",--3542
"111110001100001001000010000000000000",--3543
"111110000110000001000001100000000000",--3544
"001111001100000001000000000000000011",--3545
"111110001000001001010010000000000000",--3546
"111110000110000001000001100000000000",--3547
"001011000000000000110000000100101111",--3548
"101001000000000001010000000000000001",--3549
"000101000000000000000000111000100001",--3550
"101000000001111000000010100000000000",--3551
"000101000000000000000000111000100001",--3552
"001111001100000001100000000000000000",--3553
"011110001101000000000000000000000010",--3554
"101000000001111000000010100000000000",--3555
"000101000000000000000000111000100001",--3556
"001111001100000001110000000000000001",--3557
"111110001110001000110011100000000000",--3558
"001111001100000010000000000000000010",--3559
"111110010000001001000100000000000000",--3560
"111110001110000010000011100000000000",--3561
"001111001100000010000000000000000011",--3562
"111110010000001001010100000000000000",--3563
"111110001110000010000011100000000000",--3564
"111110000110001000110100000000000000",--3565
"001101001010000010000000000000000100",--3566
"001111010000000010010000000000000000",--3567
"111110010000001010010100000000000000",--3568
"111110001000001001000100100000000000",--3569
"001111010000000010100000000000000001",--3570
"111110010010001010100100100000000000",--3571
"111110010000000010010100000000000000",--3572
"111110001010001001010100100000000000",--3573
"001111010000000010100000000000000010",--3574
"111110010010001010100100100000000000",--3575
"111110010000000010010100000000000000",--3576
"001101001010000010000000000000000011",--3577
"011100010001000000000000000000000011",--3578
"101110010001111000000001100000000000",--3579
"011111001111000000110000000000010000",--3580
"000101000000000000000000111000001100",--3581
"111110001000001001010100100000000000",--3582
"001101001010000010000000000000001001",--3583
"001111010000000010100000000000000000",--3584
"111110010010001010100100100000000000",--3585
"111110010000000010010100000000000000",--3586
"111110001010001000110010100000000000",--3587
"001111010000000010010000000000000001",--3588
"111110001010001010010010100000000000",--3589
"111110010000000001010010100000000000",--3590
"111110000110001001000001100000000000",--3591
"001111010000000001000000000000000010",--3592
"111110000110001001000001100000000000",--3593
"111110001010000000110001100000000000",--3594
"011111001111000000110000000000000001",--3595
"111110000110010000010001100000000000",--3596
"111110001110001001110010000000000000",--3597
"111110001100001000110001100000000000",--3598
"111110001000010000110001100000000000",--3599
"010110000111000000000000000000001111",--3600
"001101001010000001010000000000000110",--3601
"011100001011000000000000000000000110",--3602
"111110000110100000000001100000000000",--3603
"111110001110010000110001100000000000",--3604
"001111001100000001000000000000000100",--3605
"111110000110001001000001100000000000",--3606
"001011000000000000110000000100101111",--3607
"000101000000000000000000111000011110",--3608
"111110000110100000000001100000000000",--3609
"111110001110000000110001100000000000",--3610
"001111001100000001000000000000000100",--3611
"111110000110001001000001100000000000",--3612
"001011000000000000110000000100101111",--3613
"101001000000000001010000000000000001",--3614
"000101000000000000000000111000100001",--3615
"101000000001111000000010100000000000",--3616
"001111000000000000110000000100101111",--3617
"010000001011000000000000000000101100",--3618
"101111001001110001001011111001001100",--3619
"101111001001100001001100110011001101",--3620
"010110001001000000110000000000101001",--3621
"001101000110000001000000000000000000",--3622
"001001111100000000111111111111111110",--3623
"010011001001000000000000000111010000",--3624
"101111001001110001000011110000100011",--3625
"101111001001100001001101011100001010",--3626
"111110000110000001000001100000000000",--3627
"001111000000000001000000000101100100",--3628
"111110001000001000110010000000000000",--3629
"001111000000000001010000000100101010",--3630
"111110001000000001010010000000000000",--3631
"001111000000000001010000000101100101",--3632
"111110001010001000110010100000000000",--3633
"001111000000000001100000000100101011",--3634
"111110001010000001100010100000000000",--3635
"001111000000000001100000000101100110",--3636
"111110001100001000110001100000000000",--3637
"001111000000000001100000000100101100",--3638
"111110000110000001100001100000000000",--3639
"001101001000000001000000000101101101",--3640
"001101001000000001010000000000000101",--3641
"001111001010000001100000000000000000",--3642
"111110001000010001100011000000000000",--3643
"001111001010000001110000000000000001",--3644
"111110001010010001110011100000000000",--3645
"001111001010000010000000000000000010",--3646
"111110000110010010000100000000000000",--3647
"001101001000000001010000000000000001",--3648
"011111001011000000010000000000011100",--3649
"101110001101111000000011000000000001",--3650
"001101001000000001010000000000000100",--3651
"001111001010000010010000000000000000",--3652
"010110010011000001100000000000010101",--3653
"101110001111111000000011000000000001",--3654
"001111001010000001110000000000000001",--3655
"010110001111000001100000000000010010",--3656
"101110010001111000000011000000000001",--3657
"001111001010000001110000000000000010",--3658
"010110001111000001100000000000001111",--3659
"001101001000000001000000000000000110",--3660
"011100001001000000000000000010100010",--3661
"000101000000000000000000111010010011",--3662
"001101001000000001000000000101101101",--3663
"001101001000000001000000000000000110",--3664
"010000001001000000000000000010100110",--3665
"101000000111111000000001000000000000",--3666
"101001000000000000010000000000000001",--3667
"001001111100000111111111111111111110",--3668
"101001111100010111100000000000000011",--3669
"000111000000000000000000100011100001",--3670
"101001111100000111100000000000000011",--3671
"001101111100000111111111111111111110",--3672
"011100000011000000000000000110011111",--3673
"000101000000000000000000111011111000",--3674
"001101001000000001000000000000000110",--3675
"011100001001000000000000000000110110",--3676
"000101000000000000000000111011110000",--3677
"011111001011000000100000000000001111",--3678
"001101001000000001010000000000000100",--3679
"001111001010000010010000000000000000",--3680
"111110010010001001100011000000000000",--3681
"001111001010000010010000000000000001",--3682
"111110010010001001110011100000000000",--3683
"111110001100000001110011000000000000",--3684
"001111001010000001110000000000000010",--3685
"111110001110001010000011100000000000",--3686
"111110001100000001110011000000000000",--3687
"001101001000000001000000000000000110",--3688
"011010001101000000000000000000000010",--3689
"011111001001000000010000000000101000",--3690
"000101000000000000000000111011110000",--3691
"011100001001000000000000000000100110",--3692
"000101000000000000000000111011110000",--3693
"111110001100001001100100100000000000",--3694
"001101001000000001100000000000000100",--3695
"001111001100000010100000000000000000",--3696
"111110010010001010100100100000000000",--3697
"111110001110001001110101000000000000",--3698
"001111001100000010110000000000000001",--3699
"111110010100001010110101000000000000",--3700
"111110010010000010100100100000000000",--3701
"111110010000001010000101000000000000",--3702
"001111001100000010110000000000000010",--3703
"111110010100001010110101000000000000",--3704
"111110010010000010100100100000000000",--3705
"001101001000000001100000000000000011",--3706
"011100001101000000000000000000000011",--3707
"101110010011111000000011000000000000",--3708
"011111001011000000110000000000010000",--3709
"000101000000000000000000111010001101",--3710
"111110001110001010000101000000000000",--3711
"001101001000000001100000000000001001",--3712
"001111001100000010110000000000000000",--3713
"111110010100001010110101000000000000",--3714
"111110010010000010100100100000000000",--3715
"111110010000001001100100000000000000",--3716
"001111001100000010100000000000000001",--3717
"111110010000001010100100000000000000",--3718
"111110010010000010000100000000000000",--3719
"111110001100001001110011000000000000",--3720
"001111001100000001110000000000000010",--3721
"111110001100001001110011000000000000",--3722
"111110010000000001100011000000000000",--3723
"011111001011000000110000000000000001",--3724
"111110001100010000010011000000000000",--3725
"001101001000000001000000000000000110",--3726
"011010001101000000000000000000000010",--3727
"011111001001000000010000000000000010",--3728
"000101000000000000000000111011110000",--3729
"010000001001000000000000000001011101",--3730
"001101000110000001000000000000000001",--3731
"010011001001000000000000000101100100",--3732
"001101001000000001000000000101101101",--3733
"001101001000000001010000000000000101",--3734
"001111001010000001100000000000000000",--3735
"111110001000010001100011000000000000",--3736
"001111001010000001110000000000000001",--3737
"111110001010010001110011100000000000",--3738
"001111001010000010000000000000000010",--3739
"111110000110010010000100000000000000",--3740
"001101001000000001010000000000000001",--3741
"011111001011000000010000000000010000",--3742
"101110001101111000000011000000000001",--3743
"001101001000000001010000000000000100",--3744
"001111001010000010010000000000000000",--3745
"010110010011000001100000000000001001",--3746
"101110001111111000000011000000000001",--3747
"001111001010000001110000000000000001",--3748
"010110001111000001100000000000000110",--3749
"101110010001111000000011000000000001",--3750
"001111001010000001110000000000000010",--3751
"010110001111000001100000000000000011",--3752
"001101001000000001000000000000000110",--3753
"011100001001000000000000000001000101",--3754
"000101000000000000000000111011100100",--3755
"001101001000000001000000000000000110",--3756
"011100001001000000000000000000110110",--3757
"000101000000000000000000111011110000",--3758
"011111001011000000100000000000001111",--3759
"001101001000000001010000000000000100",--3760
"001111001010000010010000000000000000",--3761
"111110010010001001100011000000000000",--3762
"001111001010000010010000000000000001",--3763
"111110010010001001110011100000000000",--3764
"111110001100000001110011000000000000",--3765
"001111001010000001110000000000000010",--3766
"111110001110001010000011100000000000",--3767
"111110001100000001110011000000000000",--3768
"001101001000000001000000000000000110",--3769
"011010001101000000000000000000000010",--3770
"011111001001000000010000000000101000",--3771
"000101000000000000000000111011110000",--3772
"011100001001000000000000000000100110",--3773
"000101000000000000000000111011110000",--3774
"111110001100001001100100100000000000",--3775
"001101001000000001100000000000000100",--3776
"001111001100000010100000000000000000",--3777
"111110010010001010100100100000000000",--3778
"111110001110001001110101000000000000",--3779
"001111001100000010110000000000000001",--3780
"111110010100001010110101000000000000",--3781
"111110010010000010100100100000000000",--3782
"111110010000001010000101000000000000",--3783
"001111001100000010110000000000000010",--3784
"111110010100001010110101000000000000",--3785
"111110010010000010100100100000000000",--3786
"001101001000000001100000000000000011",--3787
"011100001101000000000000000000000011",--3788
"101110010011111000000011000000000000",--3789
"011111001011000000110000000000010000",--3790
"000101000000000000000000111011011110",--3791
"111110001110001010000101000000000000",--3792
"001101001000000001100000000000001001",--3793
"001111001100000010110000000000000000",--3794
"111110010100001010110101000000000000",--3795
"111110010010000010100100100000000000",--3796
"111110010000001001100100000000000000",--3797
"001111001100000010100000000000000001",--3798
"111110010000001010100100000000000000",--3799
"111110010010000010000100000000000000",--3800
"111110001100001001110011000000000000",--3801
"001111001100000001110000000000000010",--3802
"111110001100001001110011000000000000",--3803
"111110010000000001100011000000000000",--3804
"011111001011000000110000000000000001",--3805
"111110001100010000010011000000000000",--3806
"001101001000000001000000000000000110",--3807
"011010001101000000000000000000000010",--3808
"011111001001000000010000000000000010",--3809
"000101000000000000000000111011110000",--3810
"010000001001000000000000000000001100",--3811
"101000000111111000000001000000000000",--3812
"101001000000000000010000000000000010",--3813
"101110001011111000001111100000000000",--3814
"101110000111111000000010100000000000",--3815
"101110001001111000000001100000000000",--3816
"101110111111111000000010000000000000",--3817
"001001111100000111111111111111111101",--3818
"101001111100010111100000000000000100",--3819
"000111000000000000000000011110001000",--3820
"101001111100000111100000000000000100",--3821
"001101111100000111111111111111111101",--3822
"011100000011000000000000000100001001",--3823
"101001000000000000010000000000000001",--3824
"001101111100000000101111111111111110",--3825
"001001111100000111111111111111111101",--3826
"101001111100010111100000000000000100",--3827
"000111000000000000000000100011100001",--3828
"101001111100000111100000000000000100",--3829
"001101111100000111111111111111111101",--3830
"011100000011000000000000000100000001",--3831
"001101111100000000011111111111111111",--3832
"101001000010000000010000000000000001",--3833
"001101111100000000110000000000000000",--3834
"001100000110000000010001000000000000",--3835
"011111000101000000000000000000000010",--3836
"101000000001111000000000100000000000",--3837
"000100000000000000001111100000000000",--3838
"001101000100000000100000000100110001",--3839
"001001111100000000011111111111111110",--3840
"101000000001111000000000100000000000",--3841
"001001111100000111111111111111111101",--3842
"101001111100010111100000000000000100",--3843
"000111000000000000000000100011100001",--3844
"101001111100000111100000000000000100",--3845
"001101111100000111111111111111111101",--3846
"011100000011000000000000000011101111",--3847
"001101111100000000011111111111111110",--3848
"101001000010000000010000000000000001",--3849
"001101111100000000110000000000000000",--3850
"001100000110000000010001000000000000",--3851
"011111000101000000000000000000000010",--3852
"101000000001111000000000100000000000",--3853
"000100000000000000001111100000000000",--3854
"001101000100000000100000000100110001",--3855
"001101000100000001000000000000000000",--3856
"001001111100000000011111111111111101",--3857
"010011001001000000000000000011001100",--3858
"001101001000000001010000000101101101",--3859
"001111000000000000110000000100101010",--3860
"001101001010000001100000000000000101",--3861
"001111001100000001000000000000000000",--3862
"111110000110010001000001100000000000",--3863
"001111000000000001000000000100101011",--3864
"001111001100000001010000000000000001",--3865
"111110001000010001010010000000000000",--3866
"001111000000000001010000000100101100",--3867
"001111001100000001100000000000000010",--3868
"111110001010010001100010100000000000",--3869
"001101001000000001100000000010111110",--3870
"001101001010000001110000000000000001",--3871
"011111001111000000010000000000111100",--3872
"001111001100000001100000000000000000",--3873
"111110001100010000110011000000000000",--3874
"001111001100000001110000000000000001",--3875
"111110001100001001110011000000000000",--3876
"001111000000000001110000000011111011",--3877
"111110001100001001110011100000000000",--3878
"111110001110000001000011100000000001",--3879
"001101001010000001010000000000000100",--3880
"001111001010000010000000000000000001",--3881
"010110010001000001110000000000000111",--3882
"001111000000000001110000000011111100",--3883
"111110001100001001110011100000000000",--3884
"111110001110000001010011100000000001",--3885
"001111001010000010000000000000000010",--3886
"010110010001000001110000000000000010",--3887
"001111001100000001110000000000000001",--3888
"011110001111000000000000000000101000",--3889
"001111001100000001100000000000000010",--3890
"111110001100010001000011000000000000",--3891
"001111001100000001110000000000000011",--3892
"111110001100001001110011000000000000",--3893
"001111000000000001110000000011111010",--3894
"111110001100001001110011100000000000",--3895
"111110001110000000110011100000000001",--3896
"001111001010000010000000000000000000",--3897
"010110010001000001110000000000000111",--3898
"001111000000000001110000000011111100",--3899
"111110001100001001110011100000000000",--3900
"111110001110000001010011100000000001",--3901
"001111001010000010000000000000000010",--3902
"010110010001000001110000000000000010",--3903
"001111001100000001110000000000000011",--3904
"011110001111000000000000000000010101",--3905
"001111001100000001100000000000000100",--3906
"111110001100010001010010100000000000",--3907
"001111001100000001100000000000000101",--3908
"111110001010001001100010100000000000",--3909
"001111000000000001100000000011111010",--3910
"111110001010001001100011000000000000",--3911
"111110001100000000110001100000000001",--3912
"001111001010000001100000000000000000",--3913
"010110001101000000110000000000000111",--3914
"001111000000000000110000000011111011",--3915
"111110001010001000110001100000000000",--3916
"111110000110000001000001100000000001",--3917
"001111001010000001000000000000000001",--3918
"010110001001000000110000000000000010",--3919
"001111001100000000110000000000000101",--3920
"011110000111000000000000000000000010",--3921
"101000000001111000000010100000000000",--3922
"000101000000000000000000111110101101",--3923
"001011000000000001010000000100101111",--3924
"101001000000000001010000000000000011",--3925
"000101000000000000000000111110101101",--3926
"001011000000000001100000000100101111",--3927
"101001000000000001010000000000000010",--3928
"000101000000000000000000111110101101",--3929
"001011000000000001100000000100101111",--3930
"101001000000000001010000000000000001",--3931
"000101000000000000000000111110101101",--3932
"011111001111000000100000000000001111",--3933
"001111001100000001100000000000000000",--3934
"011010001101000000000000000000001011",--3935
"001111001100000001100000000000000001",--3936
"111110001100001000110001100000000000",--3937
"001111001100000001100000000000000010",--3938
"111110001100001001000010000000000000",--3939
"111110000110000001000001100000000000",--3940
"001111001100000001000000000000000011",--3941
"111110001000001001010010000000000000",--3942
"111110000110000001000001100000000000",--3943
"001011000000000000110000000100101111",--3944
"101001000000000001010000000000000001",--3945
"000101000000000000000000111110101101",--3946
"101000000001111000000010100000000000",--3947
"000101000000000000000000111110101101",--3948
"001111001100000001100000000000000000",--3949
"011110001101000000000000000000000010",--3950
"101000000001111000000010100000000000",--3951
"000101000000000000000000111110101101",--3952
"001111001100000001110000000000000001",--3953
"111110001110001000110011100000000000",--3954
"001111001100000010000000000000000010",--3955
"111110010000001001000100000000000000",--3956
"111110001110000010000011100000000000",--3957
"001111001100000010000000000000000011",--3958
"111110010000001001010100000000000000",--3959
"111110001110000010000011100000000000",--3960
"111110000110001000110100000000000000",--3961
"001101001010000010000000000000000100",--3962
"001111010000000010010000000000000000",--3963
"111110010000001010010100000000000000",--3964
"111110001000001001000100100000000000",--3965
"001111010000000010100000000000000001",--3966
"111110010010001010100100100000000000",--3967
"111110010000000010010100000000000000",--3968
"111110001010001001010100100000000000",--3969
"001111010000000010100000000000000010",--3970
"111110010010001010100100100000000000",--3971
"111110010000000010010100000000000000",--3972
"001101001010000010000000000000000011",--3973
"011100010001000000000000000000000011",--3974
"101110010001111000000001100000000000",--3975
"011111001111000000110000000000010000",--3976
"000101000000000000000000111110011000",--3977
"111110001000001001010100100000000000",--3978
"001101001010000010000000000000001001",--3979
"001111010000000010100000000000000000",--3980
"111110010010001010100100100000000000",--3981
"111110010000000010010100000000000000",--3982
"111110001010001000110010100000000000",--3983
"001111010000000010010000000000000001",--3984
"111110001010001010010010100000000000",--3985
"111110010000000001010010100000000000",--3986
"111110000110001001000001100000000000",--3987
"001111010000000001000000000000000010",--3988
"111110000110001001000001100000000000",--3989
"111110001010000000110001100000000000",--3990
"011111001111000000110000000000000001",--3991
"111110000110010000010001100000000000",--3992
"111110001110001001110010000000000000",--3993
"111110001100001000110001100000000000",--3994
"111110001000010000110001100000000000",--3995
"010110000111000000000000000000001111",--3996
"001101001010000001010000000000000110",--3997
"011100001011000000000000000000000110",--3998
"111110000110100000000001100000000000",--3999
"111110001110010000110001100000000000",--4000
"001111001100000001000000000000000100",--4001
"111110000110001001000001100000000000",--4002
"001011000000000000110000000100101111",--4003
"000101000000000000000000111110101010",--4004
"111110000110100000000001100000000000",--4005
"111110001110000000110001100000000000",--4006
"001111001100000001000000000000000100",--4007
"111110000110001001000001100000000000",--4008
"001011000000000000110000000100101111",--4009
"101001000000000001010000000000000001",--4010
"000101000000000000000000111110101101",--4011
"101000000001111000000010100000000000",--4012
"001111000000000000110000000100101111",--4013
"010000001011000000000000000000100110",--4014
"101111001001110001001011111001001100",--4015
"101111001001100001001100110011001101",--4016
"010110001001000000110000000000100011",--4017
"101111001001110001000011110000100011",--4018
"101111001001100001001101011100001010",--4019
"111110000110000001000001100000000000",--4020
"001111000000000001000000000101100100",--4021
"111110001000001000110010000000000000",--4022
"001111000000000001010000000100101010",--4023
"111110001000000001010010000000000000",--4024
"001111000000000001010000000101100101",--4025
"111110001010001000110010100000000000",--4026
"001111000000000001100000000100101011",--4027
"111110001010000001100010100000000000",--4028
"001111000000000001100000000101100110",--4029
"111110001100001000110001100000000000",--4030
"001111000000000001100000000100101100",--4031
"111110000110000001100001100000000000",--4032
"001001111100000000101111111111111100",--4033
"101000000001111000000000100000000000",--4034
"101110001011111000001111100000000000",--4035
"101110000111111000000010100000000000",--4036
"101110001001111000000001100000000000",--4037
"101110111111111000000010000000000000",--4038
"001001111100000111111111111111111011",--4039
"101001111100010111100000000000000110",--4040
"000111000000000000000000011110001000",--4041
"101001111100000111100000000000000110",--4042
"001101111100000111111111111111111011",--4043
"011100000011000000000000000000101000",--4044
"101001000000000000010000000000000001",--4045
"001101111100000000101111111111111100",--4046
"101001111100010111100000000000000110",--4047
"000111000000000000000000100011100001",--4048
"101001111100000111100000000000000110",--4049
"001101111100000111111111111111111011",--4050
"011100000011000000000000000000100001",--4051
"000101000000000000000000111111011111",--4052
"001101001000000001000000000101101101",--4053
"001101001000000001000000000000000110",--4054
"010000001001000000000000000000000111",--4055
"101001000000000000010000000000000001",--4056
"001001111100000111111111111111111100",--4057
"101001111100010111100000000000000101",--4058
"000111000000000000000000100011100001",--4059
"101001111100000111100000000000000101",--4060
"001101111100000111111111111111111100",--4061
"011100000011000000000000000000010110",--4062
"001101111100000000011111111111111101",--4063
"101001000010000000010000000000000001",--4064
"001101111100000000110000000000000000",--4065
"001100000110000000010001000000000000",--4066
"011111000101000000000000000000000010",--4067
"101000000001111000000000100000000000",--4068
"000100000000000000001111100000000000",--4069
"001101000100000000100000000100110001",--4070
"001001111100000000011111111111111100",--4071
"101000000001111000000000100000000000",--4072
"001001111100000111111111111111111011",--4073
"101001111100010111100000000000000110",--4074
"000111000000000000000000100011100001",--4075
"101001111100000111100000000000000110",--4076
"001101111100000111111111111111111011",--4077
"011100000011000000000000000000000100",--4078
"001101111100000000011111111111111100",--4079
"101001000010000000010000000000000001",--4080
"001101111100000000100000000000000000",--4081
"000101000000000000000000110101111110",--4082
"101001000000000000010000000000000001",--4083
"000100000000000000001111100000000000",--4084
"101001000000000000010000000000000001",--4085
"000100000000000000001111100000000000",--4086
"101001000000000000010000000000000001",--4087
"000100000000000000001111100000000000",--4088
"101001000000000000010000000000000001",--4089
"000100000000000000001111100000000000",--4090
"001100000100000000010001100000000000",--4091
"001101000110000001000000000000000000",--4092
"011111001001000000000000000000000010",--4093
"101000000001111000000000100000000000",--4094
"000100000000000000001111100000000000",--4095
"001001111100000000110000000000000000",--4096
"001001111100000000101111111111111111",--4097
"001001111100000000011111111111111110",--4098
"010011001001011000110000001111101110",--4099
"001101001000000001010000000101101101",--4100
"001111000000000000110000000100101010",--4101
"001101001010000001100000000000000101",--4102
"001111001100000001000000000000000000",--4103
"111110000110010001000001100000000000",--4104
"001111000000000001000000000100101011",--4105
"001111001100000001010000000000000001",--4106
"111110001000010001010010000000000000",--4107
"001111000000000001010000000100101100",--4108
"001111001100000001100000000000000010",--4109
"111110001010010001100010100000000000",--4110
"001101001000000001000000000010111110",--4111
"001101001010000001100000000000000001",--4112
"011111001101000000010000000000110111",--4113
"001111001000000001100000000000000000",--4114
"111110001100010000110011000000000000",--4115
"001111001000000001110000000000000001",--4116
"111110001100001001110011000000000000",--4117
"001111000000000001110000000011111011",--4118
"111110001100001001110011100000000000",--4119
"111110001110000001000011100000000001",--4120
"001101001010000001010000000000000100",--4121
"001111001010000010000000000000000001",--4122
"010110010001000001110000000000000111",--4123
"001111000000000001110000000011111100",--4124
"111110001100001001110011100000000000",--4125
"111110001110000001010011100000000001",--4126
"001111001010000010000000000000000010",--4127
"010110010001000001110000000000000010",--4128
"001111001000000001110000000000000001",--4129
"011110001111000000000000000000100100",--4130
"001111001000000001100000000000000010",--4131
"111110001100010001000011000000000000",--4132
"001111001000000001110000000000000011",--4133
"111110001100001001110011000000000000",--4134
"001111000000000001110000000011111010",--4135
"111110001100001001110011100000000000",--4136
"111110001110000000110011100000000001",--4137
"001111001010000010000000000000000000",--4138
"010110010001000001110000000000000111",--4139
"001111000000000001110000000011111100",--4140
"111110001100001001110011100000000000",--4141
"111110001110000001010011100000000001",--4142
"001111001010000010000000000000000010",--4143
"010110010001000001110000000000000010",--4144
"001111001000000001110000000000000011",--4145
"011110001111000000000000000000010010",--4146
"001111001000000001100000000000000100",--4147
"111110001100010001010010100000000000",--4148
"001111001000000001100000000000000101",--4149
"111110001010001001100010100000000000",--4150
"001111000000000001100000000011111010",--4151
"111110001010001001100011000000000000",--4152
"111110001100000000110001100000000001",--4153
"001111001010000001100000000000000000",--4154
"010110001101000000110000000101000111",--4155
"001111000000000000110000000011111011",--4156
"111110001010001000110001100000000000",--4157
"111110000110000001000001100000000001",--4158
"001111001010000001000000000000000001",--4159
"010110001001000000110000000101000010",--4160
"001111001000000000110000000000000101",--4161
"010010000111000000000000000101000000",--4162
"001011000000000001010000000100101111",--4163
"000101000000000000000001000010010001",--4164
"001011000000000001100000000100101111",--4165
"000101000000000000000001000010010001",--4166
"001011000000000001100000000100101111",--4167
"000101000000000000000001000010010001",--4168
"011111001101000000100000000000001100",--4169
"001111001000000001100000000000000000",--4170
"011010001101000000000000000100110111",--4171
"001111001000000001100000000000000001",--4172
"111110001100001000110001100000000000",--4173
"001111001000000001100000000000000010",--4174
"111110001100001001000010000000000000",--4175
"111110000110000001000001100000000000",--4176
"001111001000000001000000000000000011",--4177
"111110001000001001010010000000000000",--4178
"111110000110000001000001100000000000",--4179
"001011000000000000110000000100101111",--4180
"000101000000000000000001000010010001",--4181
"001111001000000001100000000000000000",--4182
"010010001101000000000000000100101011",--4183
"001111001000000001110000000000000001",--4184
"111110001110001000110011100000000000",--4185
"001111001000000010000000000000000010",--4186
"111110010000001001000100000000000000",--4187
"111110001110000010000011100000000000",--4188
"001111001000000010000000000000000011",--4189
"111110010000001001010100000000000000",--4190
"111110001110000010000011100000000000",--4191
"111110000110001000110100000000000000",--4192
"001101001010000001110000000000000100",--4193
"001111001110000010010000000000000000",--4194
"111110010000001010010100000000000000",--4195
"111110001000001001000100100000000000",--4196
"001111001110000010100000000000000001",--4197
"111110010010001010100100100000000000",--4198
"111110010000000010010100000000000000",--4199
"111110001010001001010100100000000000",--4200
"001111001110000010100000000000000010",--4201
"111110010010001010100100100000000000",--4202
"111110010000000010010100000000000000",--4203
"001101001010000001110000000000000011",--4204
"011100001111000000000000000000000011",--4205
"101110010001111000000001100000000000",--4206
"011111001101000000110000000000010000",--4207
"000101000000000000000001000001111111",--4208
"111110001000001001010100100000000000",--4209
"001101001010000001110000000000001001",--4210
"001111001110000010100000000000000000",--4211
"111110010010001010100100100000000000",--4212
"111110010000000010010100000000000000",--4213
"111110001010001000110010100000000000",--4214
"001111001110000010010000000000000001",--4215
"111110001010001010010010100000000000",--4216
"111110010000000001010010100000000000",--4217
"111110000110001001000001100000000000",--4218
"001111001110000001000000000000000010",--4219
"111110000110001001000001100000000000",--4220
"111110001010000000110001100000000000",--4221
"011111001101000000110000000000000001",--4222
"111110000110010000010001100000000000",--4223
"111110001110001001110010000000000000",--4224
"111110001100001000110001100000000000",--4225
"111110001000010000110001100000000000",--4226
"010110000111000000000000000011111111",--4227
"001101001010000001010000000000000110",--4228
"011100001011000000000000000000000110",--4229
"111110000110100000000001100000000000",--4230
"111110001110010000110001100000000000",--4231
"001111001000000001000000000000000100",--4232
"111110000110001001000001100000000000",--4233
"001011000000000000110000000100101111",--4234
"000101000000000000000001000010010001",--4235
"111110000110100000000001100000000000",--4236
"111110001110000000110001100000000000",--4237
"001111001000000001000000000000000100",--4238
"111110000110001001000001100000000000",--4239
"001011000000000000110000000100101111",--4240
"001111000000000000110000000100101111",--4241
"101111001001110001001011110111001100",--4242
"101111001001100001001100110011001101",--4243
"010110001001000000110000000011101110",--4244
"001101000110000001000000000000000001",--4245
"010011001001000000000000000011101100",--4246
"001101001000000000100000000100110001",--4247
"101000000001111000000000100000000000",--4248
"001001111100000111111111111111111101",--4249
"101001111100010111100000000000000100",--4250
"000111000000000000000000100011100001",--4251
"101001111100000111100000000000000100",--4252
"001101111100000111111111111111111101",--4253
"011100000011000000000000001101010011",--4254
"001101111100000000010000000000000000",--4255
"001101000010000000100000000000000010",--4256
"010011000101000000000000000011100001",--4257
"001101000100000000100000000100110001",--4258
"001101000100000000110000000000000000",--4259
"010011000111000000000000000011001100",--4260
"001101000110000001000000000101101101",--4261
"001111000000000000110000000100101010",--4262
"001101001000000001010000000000000101",--4263
"001111001010000001000000000000000000",--4264
"111110000110010001000001100000000000",--4265
"001111000000000001000000000100101011",--4266
"001111001010000001010000000000000001",--4267
"111110001000010001010010000000000000",--4268
"001111000000000001010000000100101100",--4269
"001111001010000001100000000000000010",--4270
"111110001010010001100010100000000000",--4271
"001101000110000001010000000010111110",--4272
"001101001000000001100000000000000001",--4273
"011111001101000000010000000000111100",--4274
"001111001010000001100000000000000000",--4275
"111110001100010000110011000000000000",--4276
"001111001010000001110000000000000001",--4277
"111110001100001001110011000000000000",--4278
"001111000000000001110000000011111011",--4279
"111110001100001001110011100000000000",--4280
"111110001110000001000011100000000001",--4281
"001101001000000001000000000000000100",--4282
"001111001000000010000000000000000001",--4283
"010110010001000001110000000000000111",--4284
"001111000000000001110000000011111100",--4285
"111110001100001001110011100000000000",--4286
"111110001110000001010011100000000001",--4287
"001111001000000010000000000000000010",--4288
"010110010001000001110000000000000010",--4289
"001111001010000001110000000000000001",--4290
"011110001111000000000000000000101000",--4291
"001111001010000001100000000000000010",--4292
"111110001100010001000011000000000000",--4293
"001111001010000001110000000000000011",--4294
"111110001100001001110011000000000000",--4295
"001111000000000001110000000011111010",--4296
"111110001100001001110011100000000000",--4297
"111110001110000000110011100000000001",--4298
"001111001000000010000000000000000000",--4299
"010110010001000001110000000000000111",--4300
"001111000000000001110000000011111100",--4301
"111110001100001001110011100000000000",--4302
"111110001110000001010011100000000001",--4303
"001111001000000010000000000000000010",--4304
"010110010001000001110000000000000010",--4305
"001111001010000001110000000000000011",--4306
"011110001111000000000000000000010101",--4307
"001111001010000001100000000000000100",--4308
"111110001100010001010010100000000000",--4309
"001111001010000001100000000000000101",--4310
"111110001010001001100010100000000000",--4311
"001111000000000001100000000011111010",--4312
"111110001010001001100011000000000000",--4313
"111110001100000000110001100000000001",--4314
"001111001000000001100000000000000000",--4315
"010110001101000000110000000000000111",--4316
"001111000000000000110000000011111011",--4317
"111110001010001000110001100000000000",--4318
"111110000110000001000001100000000001",--4319
"001111001000000001000000000000000001",--4320
"010110001001000000110000000000000010",--4321
"001111001010000000110000000000000101",--4322
"011110000111000000000000000000000010",--4323
"101000000001111000000010000000000000",--4324
"000101000000000000000001000100111111",--4325
"001011000000000001010000000100101111",--4326
"101001000000000001000000000000000011",--4327
"000101000000000000000001000100111111",--4328
"001011000000000001100000000100101111",--4329
"101001000000000001000000000000000010",--4330
"000101000000000000000001000100111111",--4331
"001011000000000001100000000100101111",--4332
"101001000000000001000000000000000001",--4333
"000101000000000000000001000100111111",--4334
"011111001101000000100000000000001111",--4335
"001111001010000001100000000000000000",--4336
"011010001101000000000000000000001011",--4337
"001111001010000001100000000000000001",--4338
"111110001100001000110001100000000000",--4339
"001111001010000001100000000000000010",--4340
"111110001100001001000010000000000000",--4341
"111110000110000001000001100000000000",--4342
"001111001010000001000000000000000011",--4343
"111110001000001001010010000000000000",--4344
"111110000110000001000001100000000000",--4345
"001011000000000000110000000100101111",--4346
"101001000000000001000000000000000001",--4347
"000101000000000000000001000100111111",--4348
"101000000001111000000010000000000000",--4349
"000101000000000000000001000100111111",--4350
"001111001010000001100000000000000000",--4351
"011110001101000000000000000000000010",--4352
"101000000001111000000010000000000000",--4353
"000101000000000000000001000100111111",--4354
"001111001010000001110000000000000001",--4355
"111110001110001000110011100000000000",--4356
"001111001010000010000000000000000010",--4357
"111110010000001001000100000000000000",--4358
"111110001110000010000011100000000000",--4359
"001111001010000010000000000000000011",--4360
"111110010000001001010100000000000000",--4361
"111110001110000010000011100000000000",--4362
"111110000110001000110100000000000000",--4363
"001101001000000001110000000000000100",--4364
"001111001110000010010000000000000000",--4365
"111110010000001010010100000000000000",--4366
"111110001000001001000100100000000000",--4367
"001111001110000010100000000000000001",--4368
"111110010010001010100100100000000000",--4369
"111110010000000010010100000000000000",--4370
"111110001010001001010100100000000000",--4371
"001111001110000010100000000000000010",--4372
"111110010010001010100100100000000000",--4373
"111110010000000010010100000000000000",--4374
"001101001000000001110000000000000011",--4375
"011100001111000000000000000000000011",--4376
"101110010001111000000001100000000000",--4377
"011111001101000000110000000000010000",--4378
"000101000000000000000001000100101010",--4379
"111110001000001001010100100000000000",--4380
"001101001000000001110000000000001001",--4381
"001111001110000010100000000000000000",--4382
"111110010010001010100100100000000000",--4383
"111110010000000010010100000000000000",--4384
"111110001010001000110010100000000000",--4385
"001111001110000010010000000000000001",--4386
"111110001010001010010010100000000000",--4387
"111110010000000001010010100000000000",--4388
"111110000110001001000001100000000000",--4389
"001111001110000001000000000000000010",--4390
"111110000110001001000001100000000000",--4391
"111110001010000000110001100000000000",--4392
"011111001101000000110000000000000001",--4393
"111110000110010000010001100000000000",--4394
"111110001110001001110010000000000000",--4395
"111110001100001000110001100000000000",--4396
"111110001000010000110001100000000000",--4397
"010110000111000000000000000000001111",--4398
"001101001000000001000000000000000110",--4399
"011100001001000000000000000000000110",--4400
"111110000110100000000001100000000000",--4401
"111110001110010000110001100000000000",--4402
"001111001010000001000000000000000100",--4403
"111110000110001001000001100000000000",--4404
"001011000000000000110000000100101111",--4405
"000101000000000000000001000100111100",--4406
"111110000110100000000001100000000000",--4407
"111110001110000000110001100000000000",--4408
"001111001010000001000000000000000100",--4409
"111110000110001001000001100000000000",--4410
"001011000000000000110000000100101111",--4411
"101001000000000001000000000000000001",--4412
"000101000000000000000001000100111111",--4413
"101000000001111000000010000000000000",--4414
"001111000000000000110000000100101111",--4415
"010000001001000000000000000000100110",--4416
"101111001001110001001011111001001100",--4417
"101111001001100001001100110011001101",--4418
"010110001001000000110000000000100011",--4419
"101111001001110001000011110000100011",--4420
"101111001001100001001101011100001010",--4421
"111110000110000001000001100000000000",--4422
"001111000000000001000000000101100100",--4423
"111110001000001000110010000000000000",--4424
"001111000000000001010000000100101010",--4425
"111110001000000001010010000000000000",--4426
"001111000000000001010000000101100101",--4427
"111110001010001000110010100000000000",--4428
"001111000000000001100000000100101011",--4429
"111110001010000001100010100000000000",--4430
"001111000000000001100000000101100110",--4431
"111110001100001000110001100000000000",--4432
"001111000000000001100000000100101100",--4433
"111110000110000001100001100000000000",--4434
"001001111100000000101111111111111101",--4435
"101000000001111000000000100000000000",--4436
"101110001011111000001111100000000000",--4437
"101110000111111000000010100000000000",--4438
"101110001001111000000001100000000000",--4439
"101110111111111000000010000000000000",--4440
"001001111100000111111111111111111100",--4441
"101001111100010111100000000000000101",--4442
"000111000000000000000000011110001000",--4443
"101001111100000111100000000000000101",--4444
"001101111100000111111111111111111100",--4445
"011100000011000000000000001010010011",--4446
"101001000000000000010000000000000001",--4447
"001101111100000000101111111111111101",--4448
"101001111100010111100000000000000101",--4449
"000111000000000000000000100011100001",--4450
"101001111100000111100000000000000101",--4451
"001101111100000111111111111111111100",--4452
"011100000011000000000000001010001100",--4453
"000101000000000000000001000101110001",--4454
"001101000110000000110000000101101101",--4455
"001101000110000000110000000000000110",--4456
"010000000111000000000000000000000111",--4457
"101001000000000000010000000000000001",--4458
"001001111100000111111111111111111101",--4459
"101001111100010111100000000000000100",--4460
"000111000000000000000000100011100001",--4461
"101001111100000111100000000000000100",--4462
"001101111100000111111111111111111101",--4463
"011100000011000000000000001010000001",--4464
"001101111100000000010000000000000000",--4465
"001101000010000000100000000000000011",--4466
"010011000101000000000000000000001111",--4467
"001101000100000000100000000100110001",--4468
"101000000001111000000000100000000000",--4469
"001001111100000111111111111111111101",--4470
"101001111100010111100000000000000100",--4471
"000111000000000000000000100011100001",--4472
"101001111100000111100000000000000100",--4473
"001101111100000111111111111111111101",--4474
"011100000011000000000000001001110110",--4475
"101001000000000000010000000000000100",--4476
"001101111100000000100000000000000000",--4477
"101001111100010111100000000000000100",--4478
"000111000000000000000000110101111110",--4479
"101001111100000111100000000000000100",--4480
"001101111100000111111111111111111101",--4481
"011100000011000000000000001001101111",--4482
"001101111100000000011111111111111110",--4483
"101001000010000000010000000000000001",--4484
"001101111100000000111111111111111111",--4485
"001100000110000000010001000000000000",--4486
"001101000100000001000000000000000000",--4487
"011111001001000000000000000000000010",--4488
"101000000001111000000000100000000000",--4489
"000100000000000000001111100000000000",--4490
"001001111100000000101111111111111101",--4491
"001001111100000000011111111111111100",--4492
"010011001001011000110000000101111010",--4493
"001101001000000001010000000101101101",--4494
"001111000000000000110000000100101010",--4495
"001101001010000001100000000000000101",--4496
"001111001100000001000000000000000000",--4497
"111110000110010001000001100000000000",--4498
"001111000000000001000000000100101011",--4499
"001111001100000001010000000000000001",--4500
"111110001000010001010010000000000000",--4501
"001111000000000001010000000100101100",--4502
"001111001100000001100000000000000010",--4503
"111110001010010001100010100000000000",--4504
"001101001000000001000000000010111110",--4505
"001101001010000001100000000000000001",--4506
"011111001101000000010000000000110111",--4507
"001111001000000001100000000000000000",--4508
"111110001100010000110011000000000000",--4509
"001111001000000001110000000000000001",--4510
"111110001100001001110011000000000000",--4511
"001111000000000001110000000011111011",--4512
"111110001100001001110011100000000000",--4513
"111110001110000001000011100000000001",--4514
"001101001010000001010000000000000100",--4515
"001111001010000010000000000000000001",--4516
"010110010001000001110000000000000111",--4517
"001111000000000001110000000011111100",--4518
"111110001100001001110011100000000000",--4519
"111110001110000001010011100000000001",--4520
"001111001010000010000000000000000010",--4521
"010110010001000001110000000000000010",--4522
"001111001000000001110000000000000001",--4523
"011110001111000000000000000000100100",--4524
"001111001000000001100000000000000010",--4525
"111110001100010001000011000000000000",--4526
"001111001000000001110000000000000011",--4527
"111110001100001001110011000000000000",--4528
"001111000000000001110000000011111010",--4529
"111110001100001001110011100000000000",--4530
"111110001110000000110011100000000001",--4531
"001111001010000010000000000000000000",--4532
"010110010001000001110000000000000111",--4533
"001111000000000001110000000011111100",--4534
"111110001100001001110011100000000000",--4535
"111110001110000001010011100000000001",--4536
"001111001010000010000000000000000010",--4537
"010110010001000001110000000000000010",--4538
"001111001000000001110000000000000011",--4539
"011110001111000000000000000000010010",--4540
"001111001000000001100000000000000100",--4541
"111110001100010001010010100000000000",--4542
"001111001000000001100000000000000101",--4543
"111110001010001001100010100000000000",--4544
"001111000000000001100000000011111010",--4545
"111110001010001001100011000000000000",--4546
"111110001100000000110001100000000001",--4547
"001111001010000001100000000000000000",--4548
"010110001101000000110000000100111110",--4549
"001111000000000000110000000011111011",--4550
"111110001010001000110001100000000000",--4551
"111110000110000001000001100000000001",--4552
"001111001010000001000000000000000001",--4553
"010110001001000000110000000100111001",--4554
"001111001000000000110000000000000101",--4555
"010010000111000000000000000100110111",--4556
"001011000000000001010000000100101111",--4557
"000101000000000000000001001000011011",--4558
"001011000000000001100000000100101111",--4559
"000101000000000000000001001000011011",--4560
"001011000000000001100000000100101111",--4561
"000101000000000000000001001000011011",--4562
"011111001101000000100000000000001100",--4563
"001111001000000001100000000000000000",--4564
"011010001101000000000000000100101110",--4565
"001111001000000001100000000000000001",--4566
"111110001100001000110001100000000000",--4567
"001111001000000001100000000000000010",--4568
"111110001100001001000010000000000000",--4569
"111110000110000001000001100000000000",--4570
"001111001000000001000000000000000011",--4571
"111110001000001001010010000000000000",--4572
"111110000110000001000001100000000000",--4573
"001011000000000000110000000100101111",--4574
"000101000000000000000001001000011011",--4575
"001111001000000001100000000000000000",--4576
"010010001101000000000000000100100010",--4577
"001111001000000001110000000000000001",--4578
"111110001110001000110011100000000000",--4579
"001111001000000010000000000000000010",--4580
"111110010000001001000100000000000000",--4581
"111110001110000010000011100000000000",--4582
"001111001000000010000000000000000011",--4583
"111110010000001001010100000000000000",--4584
"111110001110000010000011100000000000",--4585
"111110000110001000110100000000000000",--4586
"001101001010000001110000000000000100",--4587
"001111001110000010010000000000000000",--4588
"111110010000001010010100000000000000",--4589
"111110001000001001000100100000000000",--4590
"001111001110000010100000000000000001",--4591
"111110010010001010100100100000000000",--4592
"111110010000000010010100000000000000",--4593
"111110001010001001010100100000000000",--4594
"001111001110000010100000000000000010",--4595
"111110010010001010100100100000000000",--4596
"111110010000000010010100000000000000",--4597
"001101001010000001110000000000000011",--4598
"011100001111000000000000000000000011",--4599
"101110010001111000000001100000000000",--4600
"011111001101000000110000000000010000",--4601
"000101000000000000000001001000001001",--4602
"111110001000001001010100100000000000",--4603
"001101001010000001110000000000001001",--4604
"001111001110000010100000000000000000",--4605
"111110010010001010100100100000000000",--4606
"111110010000000010010100000000000000",--4607
"111110001010001000110010100000000000",--4608
"001111001110000010010000000000000001",--4609
"111110001010001010010010100000000000",--4610
"111110010000000001010010100000000000",--4611
"111110000110001001000001100000000000",--4612
"001111001110000001000000000000000010",--4613
"111110000110001001000001100000000000",--4614
"111110001010000000110001100000000000",--4615
"011111001101000000110000000000000001",--4616
"111110000110010000010001100000000000",--4617
"111110001110001001110010000000000000",--4618
"111110001100001000110001100000000000",--4619
"111110001000010000110001100000000000",--4620
"010110000111000000000000000011110110",--4621
"001101001010000001010000000000000110",--4622
"011100001011000000000000000000000110",--4623
"111110000110100000000001100000000000",--4624
"111110001110010000110001100000000000",--4625
"001111001000000001000000000000000100",--4626
"111110000110001001000001100000000000",--4627
"001011000000000000110000000100101111",--4628
"000101000000000000000001001000011011",--4629
"111110000110100000000001100000000000",--4630
"111110001110000000110001100000000000",--4631
"001111001000000001000000000000000100",--4632
"111110000110001001000001100000000000",--4633
"001011000000000000110000000100101111",--4634
"001111000000000000110000000100101111",--4635
"101111001001110001001011110111001100",--4636
"101111001001100001001100110011001101",--4637
"010110001001000000110000000011100101",--4638
"001101000100000001000000000000000001",--4639
"010011001001000000000000000011100011",--4640
"001101001000000001000000000100110001",--4641
"001101001000000001010000000000000000",--4642
"010011001011000000000000000011001110",--4643
"001101001010000001100000000101101101",--4644
"001111000000000000110000000100101010",--4645
"001101001100000001110000000000000101",--4646
"001111001110000001000000000000000000",--4647
"111110000110010001000001100000000000",--4648
"001111000000000001000000000100101011",--4649
"001111001110000001010000000000000001",--4650
"111110001000010001010010000000000000",--4651
"001111000000000001010000000100101100",--4652
"001111001110000001100000000000000010",--4653
"111110001010010001100010100000000000",--4654
"001101001010000001110000000010111110",--4655
"001101001100000010000000000000000001",--4656
"011111010001000000010000000000111100",--4657
"001111001110000001100000000000000000",--4658
"111110001100010000110011000000000000",--4659
"001111001110000001110000000000000001",--4660
"111110001100001001110011000000000000",--4661
"001111000000000001110000000011111011",--4662
"111110001100001001110011100000000000",--4663
"111110001110000001000011100000000001",--4664
"001101001100000001100000000000000100",--4665
"001111001100000010000000000000000001",--4666
"010110010001000001110000000000000111",--4667
"001111000000000001110000000011111100",--4668
"111110001100001001110011100000000000",--4669
"111110001110000001010011100000000001",--4670
"001111001100000010000000000000000010",--4671
"010110010001000001110000000000000010",--4672
"001111001110000001110000000000000001",--4673
"011110001111000000000000000000101000",--4674
"001111001110000001100000000000000010",--4675
"111110001100010001000011000000000000",--4676
"001111001110000001110000000000000011",--4677
"111110001100001001110011000000000000",--4678
"001111000000000001110000000011111010",--4679
"111110001100001001110011100000000000",--4680
"111110001110000000110011100000000001",--4681
"001111001100000010000000000000000000",--4682
"010110010001000001110000000000000111",--4683
"001111000000000001110000000011111100",--4684
"111110001100001001110011100000000000",--4685
"111110001110000001010011100000000001",--4686
"001111001100000010000000000000000010",--4687
"010110010001000001110000000000000010",--4688
"001111001110000001110000000000000011",--4689
"011110001111000000000000000000010101",--4690
"001111001110000001100000000000000100",--4691
"111110001100010001010010100000000000",--4692
"001111001110000001100000000000000101",--4693
"111110001010001001100010100000000000",--4694
"001111000000000001100000000011111010",--4695
"111110001010001001100011000000000000",--4696
"111110001100000000110001100000000001",--4697
"001111001100000001100000000000000000",--4698
"010110001101000000110000000000000111",--4699
"001111000000000000110000000011111011",--4700
"111110001010001000110001100000000000",--4701
"111110000110000001000001100000000001",--4702
"001111001100000001000000000000000001",--4703
"010110001001000000110000000000000010",--4704
"001111001110000000110000000000000101",--4705
"011110000111000000000000000000000010",--4706
"101000000001111000000011000000000000",--4707
"000101000000000000000001001010111110",--4708
"001011000000000001010000000100101111",--4709
"101001000000000001100000000000000011",--4710
"000101000000000000000001001010111110",--4711
"001011000000000001100000000100101111",--4712
"101001000000000001100000000000000010",--4713
"000101000000000000000001001010111110",--4714
"001011000000000001100000000100101111",--4715
"101001000000000001100000000000000001",--4716
"000101000000000000000001001010111110",--4717
"011111010001000000100000000000001111",--4718
"001111001110000001100000000000000000",--4719
"011010001101000000000000000000001011",--4720
"001111001110000001100000000000000001",--4721
"111110001100001000110001100000000000",--4722
"001111001110000001100000000000000010",--4723
"111110001100001001000010000000000000",--4724
"111110000110000001000001100000000000",--4725
"001111001110000001000000000000000011",--4726
"111110001000001001010010000000000000",--4727
"111110000110000001000001100000000000",--4728
"001011000000000000110000000100101111",--4729
"101001000000000001100000000000000001",--4730
"000101000000000000000001001010111110",--4731
"101000000001111000000011000000000000",--4732
"000101000000000000000001001010111110",--4733
"001111001110000001100000000000000000",--4734
"011110001101000000000000000000000010",--4735
"101000000001111000000011000000000000",--4736
"000101000000000000000001001010111110",--4737
"001111001110000001110000000000000001",--4738
"111110001110001000110011100000000000",--4739
"001111001110000010000000000000000010",--4740
"111110010000001001000100000000000000",--4741
"111110001110000010000011100000000000",--4742
"001111001110000010000000000000000011",--4743
"111110010000001001010100000000000000",--4744
"111110001110000010000011100000000000",--4745
"111110000110001000110100000000000000",--4746
"001101001100000010010000000000000100",--4747
"001111010010000010010000000000000000",--4748
"111110010000001010010100000000000000",--4749
"111110001000001001000100100000000000",--4750
"001111010010000010100000000000000001",--4751
"111110010010001010100100100000000000",--4752
"111110010000000010010100000000000000",--4753
"111110001010001001010100100000000000",--4754
"001111010010000010100000000000000010",--4755
"111110010010001010100100100000000000",--4756
"111110010000000010010100000000000000",--4757
"001101001100000010010000000000000011",--4758
"011100010011000000000000000000000011",--4759
"101110010001111000000001100000000000",--4760
"011111010001000000110000000000010000",--4761
"000101000000000000000001001010101001",--4762
"111110001000001001010100100000000000",--4763
"001101001100000010010000000000001001",--4764
"001111010010000010100000000000000000",--4765
"111110010010001010100100100000000000",--4766
"111110010000000010010100000000000000",--4767
"111110001010001000110010100000000000",--4768
"001111010010000010010000000000000001",--4769
"111110001010001010010010100000000000",--4770
"111110010000000001010010100000000000",--4771
"111110000110001001000001100000000000",--4772
"001111010010000001000000000000000010",--4773
"111110000110001001000001100000000000",--4774
"111110001010000000110001100000000000",--4775
"011111010001000000110000000000000001",--4776
"111110000110010000010001100000000000",--4777
"111110001110001001110010000000000000",--4778
"111110001100001000110001100000000000",--4779
"111110001000010000110001100000000000",--4780
"010110000111000000000000000000001111",--4781
"001101001100000001100000000000000110",--4782
"011100001101000000000000000000000110",--4783
"111110000110100000000001100000000000",--4784
"111110001110010000110001100000000000",--4785
"001111001110000001000000000000000100",--4786
"111110000110001001000001100000000000",--4787
"001011000000000000110000000100101111",--4788
"000101000000000000000001001010111011",--4789
"111110000110100000000001100000000000",--4790
"111110001110000000110001100000000000",--4791
"001111001110000001000000000000000100",--4792
"111110000110001001000001100000000000",--4793
"001011000000000000110000000100101111",--4794
"101001000000000001100000000000000001",--4795
"000101000000000000000001001010111110",--4796
"101000000001111000000011000000000000",--4797
"001111000000000000110000000100101111",--4798
"010000001101000000000000000000100111",--4799
"101111001001110001001011111001001100",--4800
"101111001001100001001100110011001101",--4801
"010110001001000000110000000000100100",--4802
"101111001001110001000011110000100011",--4803
"101111001001100001001101011100001010",--4804
"111110000110000001000001100000000000",--4805
"001111000000000001000000000101100100",--4806
"111110001000001000110010000000000000",--4807
"001111000000000001010000000100101010",--4808
"111110001000000001010010000000000000",--4809
"001111000000000001010000000101100101",--4810
"111110001010001000110010100000000000",--4811
"001111000000000001100000000100101011",--4812
"111110001010000001100010100000000000",--4813
"001111000000000001100000000101100110",--4814
"111110001100001000110001100000000000",--4815
"001111000000000001100000000100101100",--4816
"111110000110000001100001100000000000",--4817
"001001111100000001001111111111111011",--4818
"101000001001111000000001000000000000",--4819
"101000000001111000000000100000000000",--4820
"101110001011111000001111100000000000",--4821
"101110000111111000000010100000000000",--4822
"101110001001111000000001100000000000",--4823
"101110111111111000000010000000000000",--4824
"001001111100000111111111111111111010",--4825
"101001111100010111100000000000000111",--4826
"000111000000000000000000011110001000",--4827
"101001111100000111100000000000000111",--4828
"001101111100000111111111111111111010",--4829
"011100000011000000000000000000101001",--4830
"101001000000000000010000000000000001",--4831
"001101111100000000101111111111111011",--4832
"101001111100010111100000000000000111",--4833
"000111000000000000000000100011100001",--4834
"101001111100000111100000000000000111",--4835
"001101111100000111111111111111111010",--4836
"011100000011000000000000000000100010",--4837
"000101000000000000000001001011110010",--4838
"001101001010000001010000000101101101",--4839
"001101001010000001010000000000000110",--4840
"010000001011000000000000000000001000",--4841
"101000001001111000000001000000000000",--4842
"101001000000000000010000000000000001",--4843
"001001111100000111111111111111111011",--4844
"101001111100010111100000000000000110",--4845
"000111000000000000000000100011100001",--4846
"101001111100000111100000000000000110",--4847
"001101111100000111111111111111111011",--4848
"011100000011000000000000000000010110",--4849
"001101111100000000011111111111111101",--4850
"001101000010000000100000000000000010",--4851
"010011000101000000000000000000001111",--4852
"001101000100000000100000000100110001",--4853
"101000000001111000000000100000000000",--4854
"001001111100000111111111111111111011",--4855
"101001111100010111100000000000000110",--4856
"000111000000000000000000100011100001",--4857
"101001111100000111100000000000000110",--4858
"001101111100000111111111111111111011",--4859
"011100000011000000000000000000001011",--4860
"101001000000000000010000000000000011",--4861
"001101111100000000101111111111111101",--4862
"101001111100010111100000000000000110",--4863
"000111000000000000000000110101111110",--4864
"101001111100000111100000000000000110",--4865
"001101111100000111111111111111111011",--4866
"011100000011000000000000000000000100",--4867
"001101111100000000011111111111111100",--4868
"101001000010000000010000000000000001",--4869
"001101111100000000101111111111111111",--4870
"000101000000000000000000111111111011",--4871
"001101111100000000011111111111111101",--4872
"001101000010000000100000000000000001",--4873
"010011000101000000000000000011100001",--4874
"001101000100000000100000000100110001",--4875
"001101000100000000110000000000000000",--4876
"010011000111000000000000000011001100",--4877
"001101000110000001000000000101101101",--4878
"001111000000000000110000000100101010",--4879
"001101001000000001010000000000000101",--4880
"001111001010000001000000000000000000",--4881
"111110000110010001000001100000000000",--4882
"001111000000000001000000000100101011",--4883
"001111001010000001010000000000000001",--4884
"111110001000010001010010000000000000",--4885
"001111000000000001010000000100101100",--4886
"001111001010000001100000000000000010",--4887
"111110001010010001100010100000000000",--4888
"001101000110000001010000000010111110",--4889
"001101001000000001100000000000000001",--4890
"011111001101000000010000000000111100",--4891
"001111001010000001100000000000000000",--4892
"111110001100010000110011000000000000",--4893
"001111001010000001110000000000000001",--4894
"111110001100001001110011000000000000",--4895
"001111000000000001110000000011111011",--4896
"111110001100001001110011100000000000",--4897
"111110001110000001000011100000000001",--4898
"001101001000000001000000000000000100",--4899
"001111001000000010000000000000000001",--4900
"010110010001000001110000000000000111",--4901
"001111000000000001110000000011111100",--4902
"111110001100001001110011100000000000",--4903
"111110001110000001010011100000000001",--4904
"001111001000000010000000000000000010",--4905
"010110010001000001110000000000000010",--4906
"001111001010000001110000000000000001",--4907
"011110001111000000000000000000101000",--4908
"001111001010000001100000000000000010",--4909
"111110001100010001000011000000000000",--4910
"001111001010000001110000000000000011",--4911
"111110001100001001110011000000000000",--4912
"001111000000000001110000000011111010",--4913
"111110001100001001110011100000000000",--4914
"111110001110000000110011100000000001",--4915
"001111001000000010000000000000000000",--4916
"010110010001000001110000000000000111",--4917
"001111000000000001110000000011111100",--4918
"111110001100001001110011100000000000",--4919
"111110001110000001010011100000000001",--4920
"001111001000000010000000000000000010",--4921
"010110010001000001110000000000000010",--4922
"001111001010000001110000000000000011",--4923
"011110001111000000000000000000010101",--4924
"001111001010000001100000000000000100",--4925
"111110001100010001010010100000000000",--4926
"001111001010000001100000000000000101",--4927
"111110001010001001100010100000000000",--4928
"001111000000000001100000000011111010",--4929
"111110001010001001100011000000000000",--4930
"111110001100000000110001100000000001",--4931
"001111001000000001100000000000000000",--4932
"010110001101000000110000000000000111",--4933
"001111000000000000110000000011111011",--4934
"111110001010001000110001100000000000",--4935
"111110000110000001000001100000000001",--4936
"001111001000000001000000000000000001",--4937
"010110001001000000110000000000000010",--4938
"001111001010000000110000000000000101",--4939
"011110000111000000000000000000000010",--4940
"101000000001111000000010000000000000",--4941
"000101000000000000000001001110101000",--4942
"001011000000000001010000000100101111",--4943
"101001000000000001000000000000000011",--4944
"000101000000000000000001001110101000",--4945
"001011000000000001100000000100101111",--4946
"101001000000000001000000000000000010",--4947
"000101000000000000000001001110101000",--4948
"001011000000000001100000000100101111",--4949
"101001000000000001000000000000000001",--4950
"000101000000000000000001001110101000",--4951
"011111001101000000100000000000001111",--4952
"001111001010000001100000000000000000",--4953
"011010001101000000000000000000001011",--4954
"001111001010000001100000000000000001",--4955
"111110001100001000110001100000000000",--4956
"001111001010000001100000000000000010",--4957
"111110001100001001000010000000000000",--4958
"111110000110000001000001100000000000",--4959
"001111001010000001000000000000000011",--4960
"111110001000001001010010000000000000",--4961
"111110000110000001000001100000000000",--4962
"001011000000000000110000000100101111",--4963
"101001000000000001000000000000000001",--4964
"000101000000000000000001001110101000",--4965
"101000000001111000000010000000000000",--4966
"000101000000000000000001001110101000",--4967
"001111001010000001100000000000000000",--4968
"011110001101000000000000000000000010",--4969
"101000000001111000000010000000000000",--4970
"000101000000000000000001001110101000",--4971
"001111001010000001110000000000000001",--4972
"111110001110001000110011100000000000",--4973
"001111001010000010000000000000000010",--4974
"111110010000001001000100000000000000",--4975
"111110001110000010000011100000000000",--4976
"001111001010000010000000000000000011",--4977
"111110010000001001010100000000000000",--4978
"111110001110000010000011100000000000",--4979
"111110000110001000110100000000000000",--4980
"001101001000000001110000000000000100",--4981
"001111001110000010010000000000000000",--4982
"111110010000001010010100000000000000",--4983
"111110001000001001000100100000000000",--4984
"001111001110000010100000000000000001",--4985
"111110010010001010100100100000000000",--4986
"111110010000000010010100000000000000",--4987
"111110001010001001010100100000000000",--4988
"001111001110000010100000000000000010",--4989
"111110010010001010100100100000000000",--4990
"111110010000000010010100000000000000",--4991
"001101001000000001110000000000000011",--4992
"011100001111000000000000000000000011",--4993
"101110010001111000000001100000000000",--4994
"011111001101000000110000000000010000",--4995
"000101000000000000000001001110010011",--4996
"111110001000001001010100100000000000",--4997
"001101001000000001110000000000001001",--4998
"001111001110000010100000000000000000",--4999
"111110010010001010100100100000000000",--5000
"111110010000000010010100000000000000",--5001
"111110001010001000110010100000000000",--5002
"001111001110000010010000000000000001",--5003
"111110001010001010010010100000000000",--5004
"111110010000000001010010100000000000",--5005
"111110000110001001000001100000000000",--5006
"001111001110000001000000000000000010",--5007
"111110000110001001000001100000000000",--5008
"111110001010000000110001100000000000",--5009
"011111001101000000110000000000000001",--5010
"111110000110010000010001100000000000",--5011
"111110001110001001110010000000000000",--5012
"111110001100001000110001100000000000",--5013
"111110001000010000110001100000000000",--5014
"010110000111000000000000000000001111",--5015
"001101001000000001000000000000000110",--5016
"011100001001000000000000000000000110",--5017
"111110000110100000000001100000000000",--5018
"111110001110010000110001100000000000",--5019
"001111001010000001000000000000000100",--5020
"111110000110001001000001100000000000",--5021
"001011000000000000110000000100101111",--5022
"000101000000000000000001001110100101",--5023
"111110000110100000000001100000000000",--5024
"111110001110000000110001100000000000",--5025
"001111001010000001000000000000000100",--5026
"111110000110001001000001100000000000",--5027
"001011000000000000110000000100101111",--5028
"101001000000000001000000000000000001",--5029
"000101000000000000000001001110101000",--5030
"101000000001111000000010000000000000",--5031
"001111000000000000110000000100101111",--5032
"010000001001000000000000000000100110",--5033
"101111001001110001001011111001001100",--5034
"101111001001100001001100110011001101",--5035
"010110001001000000110000000000100011",--5036
"101111001001110001000011110000100011",--5037
"101111001001100001001101011100001010",--5038
"111110000110000001000001100000000000",--5039
"001111000000000001000000000101100100",--5040
"111110001000001000110010000000000000",--5041
"001111000000000001010000000100101010",--5042
"111110001000000001010010000000000000",--5043
"001111000000000001010000000101100101",--5044
"111110001010001000110010100000000000",--5045
"001111000000000001100000000100101011",--5046
"111110001010000001100010100000000000",--5047
"001111000000000001100000000101100110",--5048
"111110001100001000110001100000000000",--5049
"001111000000000001100000000100101100",--5050
"111110000110000001100001100000000000",--5051
"001001111100000000101111111111111011",--5052
"101000000001111000000000100000000000",--5053
"101110001011111000001111100000000000",--5054
"101110000111111000000010100000000000",--5055
"101110001001111000000001100000000000",--5056
"101110111111111000000010000000000000",--5057
"001001111100000111111111111111111010",--5058
"101001111100010111100000000000000111",--5059
"000111000000000000000000011110001000",--5060
"101001111100000111100000000000000111",--5061
"001101111100000111111111111111111010",--5062
"011100000011000000000000000000101000",--5063
"101001000000000000010000000000000001",--5064
"001101111100000000101111111111111011",--5065
"101001111100010111100000000000000111",--5066
"000111000000000000000000100011100001",--5067
"101001111100000111100000000000000111",--5068
"001101111100000111111111111111111010",--5069
"011100000011000000000000000000100001",--5070
"000101000000000000000001001111011010",--5071
"001101000110000000110000000101101101",--5072
"001101000110000000110000000000000110",--5073
"010000000111000000000000000000000111",--5074
"101001000000000000010000000000000001",--5075
"001001111100000111111111111111111011",--5076
"101001111100010111100000000000000110",--5077
"000111000000000000000000100011100001",--5078
"101001111100000111100000000000000110",--5079
"001101111100000111111111111111111011",--5080
"011100000011000000000000000000010110",--5081
"001101111100000000011111111111111101",--5082
"001101000010000000100000000000000010",--5083
"010011000101000000000000000000001111",--5084
"001101000100000000100000000100110001",--5085
"101000000001111000000000100000000000",--5086
"001001111100000111111111111111111011",--5087
"101001111100010111100000000000000110",--5088
"000111000000000000000000100011100001",--5089
"101001111100000111100000000000000110",--5090
"001101111100000111111111111111111011",--5091
"011100000011000000000000000000001011",--5092
"101001000000000000010000000000000011",--5093
"001101111100000000101111111111111101",--5094
"101001111100010111100000000000000110",--5095
"000111000000000000000000110101111110",--5096
"101001111100000111100000000000000110",--5097
"001101111100000111111111111111111011",--5098
"011100000011000000000000000000000100",--5099
"001101111100000000011111111111111100",--5100
"101001000010000000010000000000000001",--5101
"001101111100000000101111111111111111",--5102
"000101000000000000000000111111111011",--5103
"101001000000000000010000000000000001",--5104
"000100000000000000001111100000000000",--5105
"001101111100000000010000000000000000",--5106
"001101000010000000100000000000000001",--5107
"010011000101000000000000000011101100",--5108
"001101000100000000100000000100110001",--5109
"101000000001111000000000100000000000",--5110
"001001111100000111111111111111111101",--5111
"101001111100010111100000000000000100",--5112
"000111000000000000000000100011100001",--5113
"101001111100000111100000000000000100",--5114
"001101111100000111111111111111111101",--5115
"011100000011000000000000001101010011",--5116
"001101111100000000010000000000000000",--5117
"001101000010000000100000000000000010",--5118
"010011000101000000000000000011100001",--5119
"001101000100000000100000000100110001",--5120
"001101000100000000110000000000000000",--5121
"010011000111000000000000000011001100",--5122
"001101000110000001000000000101101101",--5123
"001111000000000000110000000100101010",--5124
"001101001000000001010000000000000101",--5125
"001111001010000001000000000000000000",--5126
"111110000110010001000001100000000000",--5127
"001111000000000001000000000100101011",--5128
"001111001010000001010000000000000001",--5129
"111110001000010001010010000000000000",--5130
"001111000000000001010000000100101100",--5131
"001111001010000001100000000000000010",--5132
"111110001010010001100010100000000000",--5133
"001101000110000001010000000010111110",--5134
"001101001000000001100000000000000001",--5135
"011111001101000000010000000000111100",--5136
"001111001010000001100000000000000000",--5137
"111110001100010000110011000000000000",--5138
"001111001010000001110000000000000001",--5139
"111110001100001001110011000000000000",--5140
"001111000000000001110000000011111011",--5141
"111110001100001001110011100000000000",--5142
"111110001110000001000011100000000001",--5143
"001101001000000001000000000000000100",--5144
"001111001000000010000000000000000001",--5145
"010110010001000001110000000000000111",--5146
"001111000000000001110000000011111100",--5147
"111110001100001001110011100000000000",--5148
"111110001110000001010011100000000001",--5149
"001111001000000010000000000000000010",--5150
"010110010001000001110000000000000010",--5151
"001111001010000001110000000000000001",--5152
"011110001111000000000000000000101000",--5153
"001111001010000001100000000000000010",--5154
"111110001100010001000011000000000000",--5155
"001111001010000001110000000000000011",--5156
"111110001100001001110011000000000000",--5157
"001111000000000001110000000011111010",--5158
"111110001100001001110011100000000000",--5159
"111110001110000000110011100000000001",--5160
"001111001000000010000000000000000000",--5161
"010110010001000001110000000000000111",--5162
"001111000000000001110000000011111100",--5163
"111110001100001001110011100000000000",--5164
"111110001110000001010011100000000001",--5165
"001111001000000010000000000000000010",--5166
"010110010001000001110000000000000010",--5167
"001111001010000001110000000000000011",--5168
"011110001111000000000000000000010101",--5169
"001111001010000001100000000000000100",--5170
"111110001100010001010010100000000000",--5171
"001111001010000001100000000000000101",--5172
"111110001010001001100010100000000000",--5173
"001111000000000001100000000011111010",--5174
"111110001010001001100011000000000000",--5175
"111110001100000000110001100000000001",--5176
"001111001000000001100000000000000000",--5177
"010110001101000000110000000000000111",--5178
"001111000000000000110000000011111011",--5179
"111110001010001000110001100000000000",--5180
"111110000110000001000001100000000001",--5181
"001111001000000001000000000000000001",--5182
"010110001001000000110000000000000010",--5183
"001111001010000000110000000000000101",--5184
"011110000111000000000000000000000010",--5185
"101000000001111000000010000000000000",--5186
"000101000000000000000001010010011101",--5187
"001011000000000001010000000100101111",--5188
"101001000000000001000000000000000011",--5189
"000101000000000000000001010010011101",--5190
"001011000000000001100000000100101111",--5191
"101001000000000001000000000000000010",--5192
"000101000000000000000001010010011101",--5193
"001011000000000001100000000100101111",--5194
"101001000000000001000000000000000001",--5195
"000101000000000000000001010010011101",--5196
"011111001101000000100000000000001111",--5197
"001111001010000001100000000000000000",--5198
"011010001101000000000000000000001011",--5199
"001111001010000001100000000000000001",--5200
"111110001100001000110001100000000000",--5201
"001111001010000001100000000000000010",--5202
"111110001100001001000010000000000000",--5203
"111110000110000001000001100000000000",--5204
"001111001010000001000000000000000011",--5205
"111110001000001001010010000000000000",--5206
"111110000110000001000001100000000000",--5207
"001011000000000000110000000100101111",--5208
"101001000000000001000000000000000001",--5209
"000101000000000000000001010010011101",--5210
"101000000001111000000010000000000000",--5211
"000101000000000000000001010010011101",--5212
"001111001010000001100000000000000000",--5213
"011110001101000000000000000000000010",--5214
"101000000001111000000010000000000000",--5215
"000101000000000000000001010010011101",--5216
"001111001010000001110000000000000001",--5217
"111110001110001000110011100000000000",--5218
"001111001010000010000000000000000010",--5219
"111110010000001001000100000000000000",--5220
"111110001110000010000011100000000000",--5221
"001111001010000010000000000000000011",--5222
"111110010000001001010100000000000000",--5223
"111110001110000010000011100000000000",--5224
"111110000110001000110100000000000000",--5225
"001101001000000001110000000000000100",--5226
"001111001110000010010000000000000000",--5227
"111110010000001010010100000000000000",--5228
"111110001000001001000100100000000000",--5229
"001111001110000010100000000000000001",--5230
"111110010010001010100100100000000000",--5231
"111110010000000010010100000000000000",--5232
"111110001010001001010100100000000000",--5233
"001111001110000010100000000000000010",--5234
"111110010010001010100100100000000000",--5235
"111110010000000010010100000000000000",--5236
"001101001000000001110000000000000011",--5237
"011100001111000000000000000000000011",--5238
"101110010001111000000001100000000000",--5239
"011111001101000000110000000000010000",--5240
"000101000000000000000001010010001000",--5241
"111110001000001001010100100000000000",--5242
"001101001000000001110000000000001001",--5243
"001111001110000010100000000000000000",--5244
"111110010010001010100100100000000000",--5245
"111110010000000010010100000000000000",--5246
"111110001010001000110010100000000000",--5247
"001111001110000010010000000000000001",--5248
"111110001010001010010010100000000000",--5249
"111110010000000001010010100000000000",--5250
"111110000110001001000001100000000000",--5251
"001111001110000001000000000000000010",--5252
"111110000110001001000001100000000000",--5253
"111110001010000000110001100000000000",--5254
"011111001101000000110000000000000001",--5255
"111110000110010000010001100000000000",--5256
"111110001110001001110010000000000000",--5257
"111110001100001000110001100000000000",--5258
"111110001000010000110001100000000000",--5259
"010110000111000000000000000000001111",--5260
"001101001000000001000000000000000110",--5261
"011100001001000000000000000000000110",--5262
"111110000110100000000001100000000000",--5263
"111110001110010000110001100000000000",--5264
"001111001010000001000000000000000100",--5265
"111110000110001001000001100000000000",--5266
"001011000000000000110000000100101111",--5267
"000101000000000000000001010010011010",--5268
"111110000110100000000001100000000000",--5269
"111110001110000000110001100000000000",--5270
"001111001010000001000000000000000100",--5271
"111110000110001001000001100000000000",--5272
"001011000000000000110000000100101111",--5273
"101001000000000001000000000000000001",--5274
"000101000000000000000001010010011101",--5275
"101000000001111000000010000000000000",--5276
"001111000000000000110000000100101111",--5277
"010000001001000000000000000000100110",--5278
"101111001001110001001011111001001100",--5279
"101111001001100001001100110011001101",--5280
"010110001001000000110000000000100011",--5281
"101111001001110001000011110000100011",--5282
"101111001001100001001101011100001010",--5283
"111110000110000001000001100000000000",--5284
"001111000000000001000000000101100100",--5285
"111110001000001000110010000000000000",--5286
"001111000000000001010000000100101010",--5287
"111110001000000001010010000000000000",--5288
"001111000000000001010000000101100101",--5289
"111110001010001000110010100000000000",--5290
"001111000000000001100000000100101011",--5291
"111110001010000001100010100000000000",--5292
"001111000000000001100000000101100110",--5293
"111110001100001000110001100000000000",--5294
"001111000000000001100000000100101100",--5295
"111110000110000001100001100000000000",--5296
"001001111100000000101111111111111101",--5297
"101000000001111000000000100000000000",--5298
"101110001011111000001111100000000000",--5299
"101110000111111000000010100000000000",--5300
"101110001001111000000001100000000000",--5301
"101110111111111000000010000000000000",--5302
"001001111100000111111111111111111100",--5303
"101001111100010111100000000000000101",--5304
"000111000000000000000000011110001000",--5305
"101001111100000111100000000000000101",--5306
"001101111100000111111111111111111100",--5307
"011100000011000000000000001010010011",--5308
"101001000000000000010000000000000001",--5309
"001101111100000000101111111111111101",--5310
"101001111100010111100000000000000101",--5311
"000111000000000000000000100011100001",--5312
"101001111100000111100000000000000101",--5313
"001101111100000111111111111111111100",--5314
"011100000011000000000000001010001100",--5315
"000101000000000000000001010011001111",--5316
"001101000110000000110000000101101101",--5317
"001101000110000000110000000000000110",--5318
"010000000111000000000000000000000111",--5319
"101001000000000000010000000000000001",--5320
"001001111100000111111111111111111101",--5321
"101001111100010111100000000000000100",--5322
"000111000000000000000000100011100001",--5323
"101001111100000111100000000000000100",--5324
"001101111100000111111111111111111101",--5325
"011100000011000000000000001010000001",--5326
"001101111100000000010000000000000000",--5327
"001101000010000000100000000000000011",--5328
"010011000101000000000000000000001111",--5329
"001101000100000000100000000100110001",--5330
"101000000001111000000000100000000000",--5331
"001001111100000111111111111111111101",--5332
"101001111100010111100000000000000100",--5333
"000111000000000000000000100011100001",--5334
"101001111100000111100000000000000100",--5335
"001101111100000111111111111111111101",--5336
"011100000011000000000000001001110110",--5337
"101001000000000000010000000000000100",--5338
"001101111100000000100000000000000000",--5339
"101001111100010111100000000000000100",--5340
"000111000000000000000000110101111110",--5341
"101001111100000111100000000000000100",--5342
"001101111100000111111111111111111101",--5343
"011100000011000000000000001001101111",--5344
"001101111100000000011111111111111110",--5345
"101001000010000000010000000000000001",--5346
"001101111100000000111111111111111111",--5347
"001100000110000000010001000000000000",--5348
"001101000100000001000000000000000000",--5349
"011111001001000000000000000000000010",--5350
"101000000001111000000000100000000000",--5351
"000100000000000000001111100000000000",--5352
"001001111100000000101111111111111101",--5353
"001001111100000000011111111111111100",--5354
"010011001001011000110000000101111010",--5355
"001101001000000001010000000101101101",--5356
"001111000000000000110000000100101010",--5357
"001101001010000001100000000000000101",--5358
"001111001100000001000000000000000000",--5359
"111110000110010001000001100000000000",--5360
"001111000000000001000000000100101011",--5361
"001111001100000001010000000000000001",--5362
"111110001000010001010010000000000000",--5363
"001111000000000001010000000100101100",--5364
"001111001100000001100000000000000010",--5365
"111110001010010001100010100000000000",--5366
"001101001000000001000000000010111110",--5367
"001101001010000001100000000000000001",--5368
"011111001101000000010000000000110111",--5369
"001111001000000001100000000000000000",--5370
"111110001100010000110011000000000000",--5371
"001111001000000001110000000000000001",--5372
"111110001100001001110011000000000000",--5373
"001111000000000001110000000011111011",--5374
"111110001100001001110011100000000000",--5375
"111110001110000001000011100000000001",--5376
"001101001010000001010000000000000100",--5377
"001111001010000010000000000000000001",--5378
"010110010001000001110000000000000111",--5379
"001111000000000001110000000011111100",--5380
"111110001100001001110011100000000000",--5381
"111110001110000001010011100000000001",--5382
"001111001010000010000000000000000010",--5383
"010110010001000001110000000000000010",--5384
"001111001000000001110000000000000001",--5385
"011110001111000000000000000000100100",--5386
"001111001000000001100000000000000010",--5387
"111110001100010001000011000000000000",--5388
"001111001000000001110000000000000011",--5389
"111110001100001001110011000000000000",--5390
"001111000000000001110000000011111010",--5391
"111110001100001001110011100000000000",--5392
"111110001110000000110011100000000001",--5393
"001111001010000010000000000000000000",--5394
"010110010001000001110000000000000111",--5395
"001111000000000001110000000011111100",--5396
"111110001100001001110011100000000000",--5397
"111110001110000001010011100000000001",--5398
"001111001010000010000000000000000010",--5399
"010110010001000001110000000000000010",--5400
"001111001000000001110000000000000011",--5401
"011110001111000000000000000000010010",--5402
"001111001000000001100000000000000100",--5403
"111110001100010001010010100000000000",--5404
"001111001000000001100000000000000101",--5405
"111110001010001001100010100000000000",--5406
"001111000000000001100000000011111010",--5407
"111110001010001001100011000000000000",--5408
"111110001100000000110001100000000001",--5409
"001111001010000001100000000000000000",--5410
"010110001101000000110000000100111110",--5411
"001111000000000000110000000011111011",--5412
"111110001010001000110001100000000000",--5413
"111110000110000001000001100000000001",--5414
"001111001010000001000000000000000001",--5415
"010110001001000000110000000100111001",--5416
"001111001000000000110000000000000101",--5417
"010010000111000000000000000100110111",--5418
"001011000000000001010000000100101111",--5419
"000101000000000000000001010101111001",--5420
"001011000000000001100000000100101111",--5421
"000101000000000000000001010101111001",--5422
"001011000000000001100000000100101111",--5423
"000101000000000000000001010101111001",--5424
"011111001101000000100000000000001100",--5425
"001111001000000001100000000000000000",--5426
"011010001101000000000000000100101110",--5427
"001111001000000001100000000000000001",--5428
"111110001100001000110001100000000000",--5429
"001111001000000001100000000000000010",--5430
"111110001100001001000010000000000000",--5431
"111110000110000001000001100000000000",--5432
"001111001000000001000000000000000011",--5433
"111110001000001001010010000000000000",--5434
"111110000110000001000001100000000000",--5435
"001011000000000000110000000100101111",--5436
"000101000000000000000001010101111001",--5437
"001111001000000001100000000000000000",--5438
"010010001101000000000000000100100010",--5439
"001111001000000001110000000000000001",--5440
"111110001110001000110011100000000000",--5441
"001111001000000010000000000000000010",--5442
"111110010000001001000100000000000000",--5443
"111110001110000010000011100000000000",--5444
"001111001000000010000000000000000011",--5445
"111110010000001001010100000000000000",--5446
"111110001110000010000011100000000000",--5447
"111110000110001000110100000000000000",--5448
"001101001010000001110000000000000100",--5449
"001111001110000010010000000000000000",--5450
"111110010000001010010100000000000000",--5451
"111110001000001001000100100000000000",--5452
"001111001110000010100000000000000001",--5453
"111110010010001010100100100000000000",--5454
"111110010000000010010100000000000000",--5455
"111110001010001001010100100000000000",--5456
"001111001110000010100000000000000010",--5457
"111110010010001010100100100000000000",--5458
"111110010000000010010100000000000000",--5459
"001101001010000001110000000000000011",--5460
"011100001111000000000000000000000011",--5461
"101110010001111000000001100000000000",--5462
"011111001101000000110000000000010000",--5463
"000101000000000000000001010101100111",--5464
"111110001000001001010100100000000000",--5465
"001101001010000001110000000000001001",--5466
"001111001110000010100000000000000000",--5467
"111110010010001010100100100000000000",--5468
"111110010000000010010100000000000000",--5469
"111110001010001000110010100000000000",--5470
"001111001110000010010000000000000001",--5471
"111110001010001010010010100000000000",--5472
"111110010000000001010010100000000000",--5473
"111110000110001001000001100000000000",--5474
"001111001110000001000000000000000010",--5475
"111110000110001001000001100000000000",--5476
"111110001010000000110001100000000000",--5477
"011111001101000000110000000000000001",--5478
"111110000110010000010001100000000000",--5479
"111110001110001001110010000000000000",--5480
"111110001100001000110001100000000000",--5481
"111110001000010000110001100000000000",--5482
"010110000111000000000000000011110110",--5483
"001101001010000001010000000000000110",--5484
"011100001011000000000000000000000110",--5485
"111110000110100000000001100000000000",--5486
"111110001110010000110001100000000000",--5487
"001111001000000001000000000000000100",--5488
"111110000110001001000001100000000000",--5489
"001011000000000000110000000100101111",--5490
"000101000000000000000001010101111001",--5491
"111110000110100000000001100000000000",--5492
"111110001110000000110001100000000000",--5493
"001111001000000001000000000000000100",--5494
"111110000110001001000001100000000000",--5495
"001011000000000000110000000100101111",--5496
"001111000000000000110000000100101111",--5497
"101111001001110001001011110111001100",--5498
"101111001001100001001100110011001101",--5499
"010110001001000000110000000011100101",--5500
"001101000100000001000000000000000001",--5501
"010011001001000000000000000011100011",--5502
"001101001000000001000000000100110001",--5503
"001101001000000001010000000000000000",--5504
"010011001011000000000000000011001110",--5505
"001101001010000001100000000101101101",--5506
"001111000000000000110000000100101010",--5507
"001101001100000001110000000000000101",--5508
"001111001110000001000000000000000000",--5509
"111110000110010001000001100000000000",--5510
"001111000000000001000000000100101011",--5511
"001111001110000001010000000000000001",--5512
"111110001000010001010010000000000000",--5513
"001111000000000001010000000100101100",--5514
"001111001110000001100000000000000010",--5515
"111110001010010001100010100000000000",--5516
"001101001010000001110000000010111110",--5517
"001101001100000010000000000000000001",--5518
"011111010001000000010000000000111100",--5519
"001111001110000001100000000000000000",--5520
"111110001100010000110011000000000000",--5521
"001111001110000001110000000000000001",--5522
"111110001100001001110011000000000000",--5523
"001111000000000001110000000011111011",--5524
"111110001100001001110011100000000000",--5525
"111110001110000001000011100000000001",--5526
"001101001100000001100000000000000100",--5527
"001111001100000010000000000000000001",--5528
"010110010001000001110000000000000111",--5529
"001111000000000001110000000011111100",--5530
"111110001100001001110011100000000000",--5531
"111110001110000001010011100000000001",--5532
"001111001100000010000000000000000010",--5533
"010110010001000001110000000000000010",--5534
"001111001110000001110000000000000001",--5535
"011110001111000000000000000000101000",--5536
"001111001110000001100000000000000010",--5537
"111110001100010001000011000000000000",--5538
"001111001110000001110000000000000011",--5539
"111110001100001001110011000000000000",--5540
"001111000000000001110000000011111010",--5541
"111110001100001001110011100000000000",--5542
"111110001110000000110011100000000001",--5543
"001111001100000010000000000000000000",--5544
"010110010001000001110000000000000111",--5545
"001111000000000001110000000011111100",--5546
"111110001100001001110011100000000000",--5547
"111110001110000001010011100000000001",--5548
"001111001100000010000000000000000010",--5549
"010110010001000001110000000000000010",--5550
"001111001110000001110000000000000011",--5551
"011110001111000000000000000000010101",--5552
"001111001110000001100000000000000100",--5553
"111110001100010001010010100000000000",--5554
"001111001110000001100000000000000101",--5555
"111110001010001001100010100000000000",--5556
"001111000000000001100000000011111010",--5557
"111110001010001001100011000000000000",--5558
"111110001100000000110001100000000001",--5559
"001111001100000001100000000000000000",--5560
"010110001101000000110000000000000111",--5561
"001111000000000000110000000011111011",--5562
"111110001010001000110001100000000000",--5563
"111110000110000001000001100000000001",--5564
"001111001100000001000000000000000001",--5565
"010110001001000000110000000000000010",--5566
"001111001110000000110000000000000101",--5567
"011110000111000000000000000000000010",--5568
"101000000001111000000011000000000000",--5569
"000101000000000000000001011000011100",--5570
"001011000000000001010000000100101111",--5571
"101001000000000001100000000000000011",--5572
"000101000000000000000001011000011100",--5573
"001011000000000001100000000100101111",--5574
"101001000000000001100000000000000010",--5575
"000101000000000000000001011000011100",--5576
"001011000000000001100000000100101111",--5577
"101001000000000001100000000000000001",--5578
"000101000000000000000001011000011100",--5579
"011111010001000000100000000000001111",--5580
"001111001110000001100000000000000000",--5581
"011010001101000000000000000000001011",--5582
"001111001110000001100000000000000001",--5583
"111110001100001000110001100000000000",--5584
"001111001110000001100000000000000010",--5585
"111110001100001001000010000000000000",--5586
"111110000110000001000001100000000000",--5587
"001111001110000001000000000000000011",--5588
"111110001000001001010010000000000000",--5589
"111110000110000001000001100000000000",--5590
"001011000000000000110000000100101111",--5591
"101001000000000001100000000000000001",--5592
"000101000000000000000001011000011100",--5593
"101000000001111000000011000000000000",--5594
"000101000000000000000001011000011100",--5595
"001111001110000001100000000000000000",--5596
"011110001101000000000000000000000010",--5597
"101000000001111000000011000000000000",--5598
"000101000000000000000001011000011100",--5599
"001111001110000001110000000000000001",--5600
"111110001110001000110011100000000000",--5601
"001111001110000010000000000000000010",--5602
"111110010000001001000100000000000000",--5603
"111110001110000010000011100000000000",--5604
"001111001110000010000000000000000011",--5605
"111110010000001001010100000000000000",--5606
"111110001110000010000011100000000000",--5607
"111110000110001000110100000000000000",--5608
"001101001100000010010000000000000100",--5609
"001111010010000010010000000000000000",--5610
"111110010000001010010100000000000000",--5611
"111110001000001001000100100000000000",--5612
"001111010010000010100000000000000001",--5613
"111110010010001010100100100000000000",--5614
"111110010000000010010100000000000000",--5615
"111110001010001001010100100000000000",--5616
"001111010010000010100000000000000010",--5617
"111110010010001010100100100000000000",--5618
"111110010000000010010100000000000000",--5619
"001101001100000010010000000000000011",--5620
"011100010011000000000000000000000011",--5621
"101110010001111000000001100000000000",--5622
"011111010001000000110000000000010000",--5623
"000101000000000000000001011000000111",--5624
"111110001000001001010100100000000000",--5625
"001101001100000010010000000000001001",--5626
"001111010010000010100000000000000000",--5627
"111110010010001010100100100000000000",--5628
"111110010000000010010100000000000000",--5629
"111110001010001000110010100000000000",--5630
"001111010010000010010000000000000001",--5631
"111110001010001010010010100000000000",--5632
"111110010000000001010010100000000000",--5633
"111110000110001001000001100000000000",--5634
"001111010010000001000000000000000010",--5635
"111110000110001001000001100000000000",--5636
"111110001010000000110001100000000000",--5637
"011111010001000000110000000000000001",--5638
"111110000110010000010001100000000000",--5639
"111110001110001001110010000000000000",--5640
"111110001100001000110001100000000000",--5641
"111110001000010000110001100000000000",--5642
"010110000111000000000000000000001111",--5643
"001101001100000001100000000000000110",--5644
"011100001101000000000000000000000110",--5645
"111110000110100000000001100000000000",--5646
"111110001110010000110001100000000000",--5647
"001111001110000001000000000000000100",--5648
"111110000110001001000001100000000000",--5649
"001011000000000000110000000100101111",--5650
"000101000000000000000001011000011001",--5651
"111110000110100000000001100000000000",--5652
"111110001110000000110001100000000000",--5653
"001111001110000001000000000000000100",--5654
"111110000110001001000001100000000000",--5655
"001011000000000000110000000100101111",--5656
"101001000000000001100000000000000001",--5657
"000101000000000000000001011000011100",--5658
"101000000001111000000011000000000000",--5659
"001111000000000000110000000100101111",--5660
"010000001101000000000000000000100111",--5661
"101111001001110001001011111001001100",--5662
"101111001001100001001100110011001101",--5663
"010110001001000000110000000000100100",--5664
"101111001001110001000011110000100011",--5665
"101111001001100001001101011100001010",--5666
"111110000110000001000001100000000000",--5667
"001111000000000001000000000101100100",--5668
"111110001000001000110010000000000000",--5669
"001111000000000001010000000100101010",--5670
"111110001000000001010010000000000000",--5671
"001111000000000001010000000101100101",--5672
"111110001010001000110010100000000000",--5673
"001111000000000001100000000100101011",--5674
"111110001010000001100010100000000000",--5675
"001111000000000001100000000101100110",--5676
"111110001100001000110001100000000000",--5677
"001111000000000001100000000100101100",--5678
"111110000110000001100001100000000000",--5679
"001001111100000001001111111111111011",--5680
"101000001001111000000001000000000000",--5681
"101000000001111000000000100000000000",--5682
"101110001011111000001111100000000000",--5683
"101110000111111000000010100000000000",--5684
"101110001001111000000001100000000000",--5685
"101110111111111000000010000000000000",--5686
"001001111100000111111111111111111010",--5687
"101001111100010111100000000000000111",--5688
"000111000000000000000000011110001000",--5689
"101001111100000111100000000000000111",--5690
"001101111100000111111111111111111010",--5691
"011100000011000000000000000000101001",--5692
"101001000000000000010000000000000001",--5693
"001101111100000000101111111111111011",--5694
"101001111100010111100000000000000111",--5695
"000111000000000000000000100011100001",--5696
"101001111100000111100000000000000111",--5697
"001101111100000111111111111111111010",--5698
"011100000011000000000000000000100010",--5699
"000101000000000000000001011001010000",--5700
"001101001010000001010000000101101101",--5701
"001101001010000001010000000000000110",--5702
"010000001011000000000000000000001000",--5703
"101000001001111000000001000000000000",--5704
"101001000000000000010000000000000001",--5705
"001001111100000111111111111111111011",--5706
"101001111100010111100000000000000110",--5707
"000111000000000000000000100011100001",--5708
"101001111100000111100000000000000110",--5709
"001101111100000111111111111111111011",--5710
"011100000011000000000000000000010110",--5711
"001101111100000000011111111111111101",--5712
"001101000010000000100000000000000010",--5713
"010011000101000000000000000000001111",--5714
"001101000100000000100000000100110001",--5715
"101000000001111000000000100000000000",--5716
"001001111100000111111111111111111011",--5717
"101001111100010111100000000000000110",--5718
"000111000000000000000000100011100001",--5719
"101001111100000111100000000000000110",--5720
"001101111100000111111111111111111011",--5721
"011100000011000000000000000000001011",--5722
"101001000000000000010000000000000011",--5723
"001101111100000000101111111111111101",--5724
"101001111100010111100000000000000110",--5725
"000111000000000000000000110101111110",--5726
"101001111100000111100000000000000110",--5727
"001101111100000111111111111111111011",--5728
"011100000011000000000000000000000100",--5729
"001101111100000000011111111111111100",--5730
"101001000010000000010000000000000001",--5731
"001101111100000000101111111111111111",--5732
"000101000000000000000000111111111011",--5733
"001101111100000000011111111111111101",--5734
"001101000010000000100000000000000001",--5735
"010011000101000000000000000011100001",--5736
"001101000100000000100000000100110001",--5737
"001101000100000000110000000000000000",--5738
"010011000111000000000000000011001100",--5739
"001101000110000001000000000101101101",--5740
"001111000000000000110000000100101010",--5741
"001101001000000001010000000000000101",--5742
"001111001010000001000000000000000000",--5743
"111110000110010001000001100000000000",--5744
"001111000000000001000000000100101011",--5745
"001111001010000001010000000000000001",--5746
"111110001000010001010010000000000000",--5747
"001111000000000001010000000100101100",--5748
"001111001010000001100000000000000010",--5749
"111110001010010001100010100000000000",--5750
"001101000110000001010000000010111110",--5751
"001101001000000001100000000000000001",--5752
"011111001101000000010000000000111100",--5753
"001111001010000001100000000000000000",--5754
"111110001100010000110011000000000000",--5755
"001111001010000001110000000000000001",--5756
"111110001100001001110011000000000000",--5757
"001111000000000001110000000011111011",--5758
"111110001100001001110011100000000000",--5759
"111110001110000001000011100000000001",--5760
"001101001000000001000000000000000100",--5761
"001111001000000010000000000000000001",--5762
"010110010001000001110000000000000111",--5763
"001111000000000001110000000011111100",--5764
"111110001100001001110011100000000000",--5765
"111110001110000001010011100000000001",--5766
"001111001000000010000000000000000010",--5767
"010110010001000001110000000000000010",--5768
"001111001010000001110000000000000001",--5769
"011110001111000000000000000000101000",--5770
"001111001010000001100000000000000010",--5771
"111110001100010001000011000000000000",--5772
"001111001010000001110000000000000011",--5773
"111110001100001001110011000000000000",--5774
"001111000000000001110000000011111010",--5775
"111110001100001001110011100000000000",--5776
"111110001110000000110011100000000001",--5777
"001111001000000010000000000000000000",--5778
"010110010001000001110000000000000111",--5779
"001111000000000001110000000011111100",--5780
"111110001100001001110011100000000000",--5781
"111110001110000001010011100000000001",--5782
"001111001000000010000000000000000010",--5783
"010110010001000001110000000000000010",--5784
"001111001010000001110000000000000011",--5785
"011110001111000000000000000000010101",--5786
"001111001010000001100000000000000100",--5787
"111110001100010001010010100000000000",--5788
"001111001010000001100000000000000101",--5789
"111110001010001001100010100000000000",--5790
"001111000000000001100000000011111010",--5791
"111110001010001001100011000000000000",--5792
"111110001100000000110001100000000001",--5793
"001111001000000001100000000000000000",--5794
"010110001101000000110000000000000111",--5795
"001111000000000000110000000011111011",--5796
"111110001010001000110001100000000000",--5797
"111110000110000001000001100000000001",--5798
"001111001000000001000000000000000001",--5799
"010110001001000000110000000000000010",--5800
"001111001010000000110000000000000101",--5801
"011110000111000000000000000000000010",--5802
"101000000001111000000010000000000000",--5803
"000101000000000000000001011100000110",--5804
"001011000000000001010000000100101111",--5805
"101001000000000001000000000000000011",--5806
"000101000000000000000001011100000110",--5807
"001011000000000001100000000100101111",--5808
"101001000000000001000000000000000010",--5809
"000101000000000000000001011100000110",--5810
"001011000000000001100000000100101111",--5811
"101001000000000001000000000000000001",--5812
"000101000000000000000001011100000110",--5813
"011111001101000000100000000000001111",--5814
"001111001010000001100000000000000000",--5815
"011010001101000000000000000000001011",--5816
"001111001010000001100000000000000001",--5817
"111110001100001000110001100000000000",--5818
"001111001010000001100000000000000010",--5819
"111110001100001001000010000000000000",--5820
"111110000110000001000001100000000000",--5821
"001111001010000001000000000000000011",--5822
"111110001000001001010010000000000000",--5823
"111110000110000001000001100000000000",--5824
"001011000000000000110000000100101111",--5825
"101001000000000001000000000000000001",--5826
"000101000000000000000001011100000110",--5827
"101000000001111000000010000000000000",--5828
"000101000000000000000001011100000110",--5829
"001111001010000001100000000000000000",--5830
"011110001101000000000000000000000010",--5831
"101000000001111000000010000000000000",--5832
"000101000000000000000001011100000110",--5833
"001111001010000001110000000000000001",--5834
"111110001110001000110011100000000000",--5835
"001111001010000010000000000000000010",--5836
"111110010000001001000100000000000000",--5837
"111110001110000010000011100000000000",--5838
"001111001010000010000000000000000011",--5839
"111110010000001001010100000000000000",--5840
"111110001110000010000011100000000000",--5841
"111110000110001000110100000000000000",--5842
"001101001000000001110000000000000100",--5843
"001111001110000010010000000000000000",--5844
"111110010000001010010100000000000000",--5845
"111110001000001001000100100000000000",--5846
"001111001110000010100000000000000001",--5847
"111110010010001010100100100000000000",--5848
"111110010000000010010100000000000000",--5849
"111110001010001001010100100000000000",--5850
"001111001110000010100000000000000010",--5851
"111110010010001010100100100000000000",--5852
"111110010000000010010100000000000000",--5853
"001101001000000001110000000000000011",--5854
"011100001111000000000000000000000011",--5855
"101110010001111000000001100000000000",--5856
"011111001101000000110000000000010000",--5857
"000101000000000000000001011011110001",--5858
"111110001000001001010100100000000000",--5859
"001101001000000001110000000000001001",--5860
"001111001110000010100000000000000000",--5861
"111110010010001010100100100000000000",--5862
"111110010000000010010100000000000000",--5863
"111110001010001000110010100000000000",--5864
"001111001110000010010000000000000001",--5865
"111110001010001010010010100000000000",--5866
"111110010000000001010010100000000000",--5867
"111110000110001001000001100000000000",--5868
"001111001110000001000000000000000010",--5869
"111110000110001001000001100000000000",--5870
"111110001010000000110001100000000000",--5871
"011111001101000000110000000000000001",--5872
"111110000110010000010001100000000000",--5873
"111110001110001001110010000000000000",--5874
"111110001100001000110001100000000000",--5875
"111110001000010000110001100000000000",--5876
"010110000111000000000000000000001111",--5877
"001101001000000001000000000000000110",--5878
"011100001001000000000000000000000110",--5879
"111110000110100000000001100000000000",--5880
"111110001110010000110001100000000000",--5881
"001111001010000001000000000000000100",--5882
"111110000110001001000001100000000000",--5883
"001011000000000000110000000100101111",--5884
"000101000000000000000001011100000011",--5885
"111110000110100000000001100000000000",--5886
"111110001110000000110001100000000000",--5887
"001111001010000001000000000000000100",--5888
"111110000110001001000001100000000000",--5889
"001011000000000000110000000100101111",--5890
"101001000000000001000000000000000001",--5891
"000101000000000000000001011100000110",--5892
"101000000001111000000010000000000000",--5893
"001111000000000000110000000100101111",--5894
"010000001001000000000000000000100110",--5895
"101111001001110001001011111001001100",--5896
"101111001001100001001100110011001101",--5897
"010110001001000000110000000000100011",--5898
"101111001001110001000011110000100011",--5899
"101111001001100001001101011100001010",--5900
"111110000110000001000001100000000000",--5901
"001111000000000001000000000101100100",--5902
"111110001000001000110010000000000000",--5903
"001111000000000001010000000100101010",--5904
"111110001000000001010010000000000000",--5905
"001111000000000001010000000101100101",--5906
"111110001010001000110010100000000000",--5907
"001111000000000001100000000100101011",--5908
"111110001010000001100010100000000000",--5909
"001111000000000001100000000101100110",--5910
"111110001100001000110001100000000000",--5911
"001111000000000001100000000100101100",--5912
"111110000110000001100001100000000000",--5913
"001001111100000000101111111111111011",--5914
"101000000001111000000000100000000000",--5915
"101110001011111000001111100000000000",--5916
"101110000111111000000010100000000000",--5917
"101110001001111000000001100000000000",--5918
"101110111111111000000010000000000000",--5919
"001001111100000111111111111111111010",--5920
"101001111100010111100000000000000111",--5921
"000111000000000000000000011110001000",--5922
"101001111100000111100000000000000111",--5923
"001101111100000111111111111111111010",--5924
"011100000011000000000000000000101000",--5925
"101001000000000000010000000000000001",--5926
"001101111100000000101111111111111011",--5927
"101001111100010111100000000000000111",--5928
"000111000000000000000000100011100001",--5929
"101001111100000111100000000000000111",--5930
"001101111100000111111111111111111010",--5931
"011100000011000000000000000000100001",--5932
"000101000000000000000001011100111000",--5933
"001101000110000000110000000101101101",--5934
"001101000110000000110000000000000110",--5935
"010000000111000000000000000000000111",--5936
"101001000000000000010000000000000001",--5937
"001001111100000111111111111111111011",--5938
"101001111100010111100000000000000110",--5939
"000111000000000000000000100011100001",--5940
"101001111100000111100000000000000110",--5941
"001101111100000111111111111111111011",--5942
"011100000011000000000000000000010110",--5943
"001101111100000000011111111111111101",--5944
"001101000010000000100000000000000010",--5945
"010011000101000000000000000000001111",--5946
"001101000100000000100000000100110001",--5947
"101000000001111000000000100000000000",--5948
"001001111100000111111111111111111011",--5949
"101001111100010111100000000000000110",--5950
"000111000000000000000000100011100001",--5951
"101001111100000111100000000000000110",--5952
"001101111100000111111111111111111011",--5953
"011100000011000000000000000000001011",--5954
"101001000000000000010000000000000011",--5955
"001101111100000000101111111111111101",--5956
"101001111100010111100000000000000110",--5957
"000111000000000000000000110101111110",--5958
"101001111100000111100000000000000110",--5959
"001101111100000111111111111111111011",--5960
"011100000011000000000000000000000100",--5961
"001101111100000000011111111111111100",--5962
"101001000010000000010000000000000001",--5963
"001101111100000000101111111111111111",--5964
"000101000000000000000000111111111011",--5965
"101001000000000000010000000000000001",--5966
"000100000000000000001111100000000000",--5967
"101001000000000000010000000000000001",--5968
"000100000000000000001111100000000000",--5969
"001100000100000000010010000000000000",--5970
"010011001000000000001111100000000000",--5971
"001101001000000001010000000101101101",--5972
"001111000000000000110000000100010101",--5973
"001101001010000001100000000000000101",--5974
"001111001100000001000000000000000000",--5975
"111110000110010001000001100000000000",--5976
"001111000000000001000000000100010110",--5977
"001111001100000001010000000000000001",--5978
"111110001000010001010010000000000000",--5979
"001111000000000001010000000100010111",--5980
"001111001100000001100000000000000010",--5981
"111110001010010001100010100000000000",--5982
"001101001010000001100000000000000001",--5983
"011111001101000000010000000001010100",--5984
"001111000110000001100000000000000000",--5985
"010010001101000000000000000000011010",--5986
"001101001010000001100000000000000100",--5987
"001101001010000001110000000000000110",--5988
"011010001101000000000000000000000010",--5989
"101001000000000010000000000000000001",--5990
"000101000000000000000001011101101001",--5991
"101000000001111000000100000000000000",--5992
"001111001100000001100000000000000000",--5993
"011100001111000010000000000000000001",--5994
"101110001101111000000011000000000010",--5995
"111110001100010000110011000000000000",--5996
"001111000110000001110000000000000000",--5997
"111110001110011000000011100000000000",--5998
"111110001100001001110011000000000000",--5999
"001111000110000001110000000000000001",--6000
"111110001100001001110011100000000000",--6001
"111110001110000001000011100000000001",--6002
"001111001100000010000000000000000001",--6003
"010110010001000001110000000000001000",--6004
"001111000110000001110000000000000010",--6005
"111110001100001001110011100000000000",--6006
"111110001110000001010011100000000001",--6007
"001111001100000010000000000000000010",--6008
"010110010001000001110000000000000011",--6009
"001011000000000001100000000100101111",--6010
"101001000000000001010000000000000001",--6011
"000101000000000000000001101000011000",--6012
"001111000110000001100000000000000001",--6013
"010010001101000000000000000000011010",--6014
"001101001010000001100000000000000100",--6015
"001101001010000001110000000000000110",--6016
"011010001101000000000000000000000010",--6017
"101001000000000010000000000000000001",--6018
"000101000000000000000001011110000101",--6019
"101000000001111000000100000000000000",--6020
"001111001100000001100000000000000001",--6021
"011100001111000010000000000000000001",--6022
"101110001101111000000011000000000010",--6023
"111110001100010001000011000000000000",--6024
"001111000110000001110000000000000001",--6025
"111110001110011000000011100000000000",--6026
"111110001100001001110011000000000000",--6027
"001111000110000001110000000000000010",--6028
"111110001100001001110011100000000000",--6029
"111110001110000001010011100000000001",--6030
"001111001100000010000000000000000010",--6031
"010110010001000001110000000000001000",--6032
"001111000110000001110000000000000000",--6033
"111110001100001001110011100000000000",--6034
"111110001110000000110011100000000001",--6035
"001111001100000010000000000000000000",--6036
"010110010001000001110000000000000011",--6037
"001011000000000001100000000100101111",--6038
"101001000000000001010000000000000010",--6039
"000101000000000000000001101000011000",--6040
"001111000110000001100000000000000010",--6041
"010010001101000000000000000010101001",--6042
"001101001010000001100000000000000100",--6043
"001101001010000001010000000000000110",--6044
"011010001101000000000000000000000010",--6045
"101001000000000001110000000000000001",--6046
"000101000000000000000001011110100001",--6047
"101000000001111000000011100000000000",--6048
"001111001100000001100000000000000010",--6049
"011100001011000001110000000000000001",--6050
"101110001101111000000011000000000010",--6051
"111110001100010001010010100000000000",--6052
"001111000110000001100000000000000010",--6053
"111110001100011000000011000000000000",--6054
"111110001010001001100010100000000000",--6055
"001111000110000001100000000000000000",--6056
"111110001010001001100011000000000000",--6057
"111110001100000000110001100000000001",--6058
"001111001100000001100000000000000000",--6059
"010110001101000000110000000010010111",--6060
"001111000110000000110000000000000001",--6061
"111110001010001000110001100000000000",--6062
"111110000110000001000001100000000001",--6063
"001111001100000001000000000000000001",--6064
"010110001001000000110000000010010010",--6065
"001011000000000001010000000100101111",--6066
"101001000000000001010000000000000011",--6067
"000101000000000000000001101000011000",--6068
"011111001101000000100000000000011010",--6069
"001101001010000001010000000000000100",--6070
"001111000110000001100000000000000000",--6071
"001111001010000001110000000000000000",--6072
"111110001100001001110011000000000000",--6073
"001111000110000001110000000000000001",--6074
"001111001010000010000000000000000001",--6075
"111110001110001010000011100000000000",--6076
"111110001100000001110011000000000000",--6077
"001111000110000001110000000000000010",--6078
"001111001010000010000000000000000010",--6079
"111110001110001010000011100000000000",--6080
"111110001100000001110011000000000000",--6081
"010110001101000000000000000010000001",--6082
"001111001010000001110000000000000000",--6083
"111110001110001000110001100000000000",--6084
"001111001010000001110000000000000001",--6085
"111110001110001001000010000000000000",--6086
"111110000110000001000001100000000000",--6087
"001111001010000001000000000000000010",--6088
"111110001000001001010010000000000000",--6089
"111110000110000001000001100000000010",--6090
"111110001100011000000010000000000000",--6091
"111110000110001001000001100000000000",--6092
"001011000000000000110000000100101111",--6093
"101001000000000001010000000000000001",--6094
"000101000000000000000001101000011000",--6095
"001111000110000001100000000000000000",--6096
"001111000110000001110000000000000001",--6097
"001111000110000010000000000000000010",--6098
"111110001100001001100100100000000000",--6099
"001101001010000001110000000000000100",--6100
"001111001110000010100000000000000000",--6101
"111110010010001010100100100000000000",--6102
"111110001110001001110101000000000000",--6103
"001111001110000010110000000000000001",--6104
"111110010100001010110101000000000000",--6105
"111110010010000010100100100000000000",--6106
"111110010000001010000101000000000000",--6107
"001111001110000010110000000000000010",--6108
"111110010100001010110101000000000000",--6109
"111110010010000010100100100000000000",--6110
"001101001010000010000000000000000011",--6111
"011100010001000000000000000000000011",--6112
"101110010011111000000011000000000000",--6113
"011110010011000000000000000000001111",--6114
"000101000000000000000001100001000100",--6115
"111110001110001010000101000000000000",--6116
"001101001010000010010000000000001001",--6117
"001111010010000010110000000000000000",--6118
"111110010100001010110101000000000000",--6119
"111110010010000010100100100000000000",--6120
"111110010000001001100100000000000000",--6121
"001111010010000010100000000000000001",--6122
"111110010000001010100100000000000000",--6123
"111110010010000010000100000000000000",--6124
"111110001100001001110011000000000000",--6125
"001111010010000001110000000000000010",--6126
"111110001100001001110011000000000000",--6127
"111110010000000001100011000000000000",--6128
"010010001101000000000000000001010010",--6129
"001111000110000001110000000000000000",--6130
"001111000110000010000000000000000001",--6131
"001111000110000010010000000000000010",--6132
"111110001110001000110101000000000000",--6133
"001111001110000010110000000000000000",--6134
"111110010100001010110101000000000000",--6135
"111110010000001001000101100000000000",--6136
"001111001110000011000000000000000001",--6137
"111110010110001011000101100000000000",--6138
"111110010100000010110101000000000000",--6139
"111110010010001001010101100000000000",--6140
"001111001110000011000000000000000010",--6141
"111110010110001011000101100000000000",--6142
"111110010100000010110101000000000000",--6143
"011100010001000000000000000000000010",--6144
"101110010101111000000011100000000000",--6145
"000101000000000000000001100000011000",--6146
"111110010010001001000101100000000000",--6147
"111110010000001001010110000000000000",--6148
"111110010110000011000101100000000000",--6149
"001101001010000010010000000000001001",--6150
"001111010010000011000000000000000000",--6151
"111110010110001011000101100000000000",--6152
"111110001110001001010110000000000000",--6153
"111110010010001000110100100000000000",--6154
"111110011000000010010100100000000000",--6155
"001111010010000011000000000000000001",--6156
"111110010010001011000100100000000000",--6157
"111110010110000010010100100000000000",--6158
"111110001110001001000011100000000000",--6159
"111110010000001000110100000000000000",--6160
"111110001110000010000011100000000000",--6161
"001111010010000010000000000000000010",--6162
"111110001110001010000011100000000000",--6163
"111110010010000001110011100000000000",--6164
"101111000001110010000011111100000000",--6165
"111110001110001010000011100000000000",--6166
"111110010100000001110011100000000000",--6167
"111110000110001000110100000000000000",--6168
"001111001110000010010000000000000000",--6169
"111110010000001010010100000000000000",--6170
"111110001000001001000100100000000000",--6171
"001111001110000010100000000000000001",--6172
"111110010010001010100100100000000000",--6173
"111110010000000010010100000000000000",--6174
"111110001010001001010100100000000000",--6175
"001111001110000010100000000000000010",--6176
"111110010010001010100100100000000000",--6177
"111110010000000010010100000000000000",--6178
"011100010001000000000000000000000011",--6179
"101110010001111000000001100000000000",--6180
"011111001101000000110000000000010000",--6181
"000101000000000000000001100000110101",--6182
"111110001000001001010100100000000000",--6183
"001101001010000001110000000000001001",--6184
"001111001110000010100000000000000000",--6185
"111110010010001010100100100000000000",--6186
"111110010000000010010100000000000000",--6187
"111110001010001000110010100000000000",--6188
"001111001110000010010000000000000001",--6189
"111110001010001010010010100000000000",--6190
"111110010000000001010010100000000000",--6191
"111110000110001001000001100000000000",--6192
"001111001110000001000000000000000010",--6193
"111110000110001001000001100000000000",--6194
"111110001010000000110001100000000000",--6195
"011111001101000000110000000000000001",--6196
"111110000110010000010001100000000000",--6197
"111110001110001001110010000000000000",--6198
"111110001100001000110001100000000000",--6199
"111110001000010000110001100000000000",--6200
"010110000111000000000000000000001010",--6201
"111110000110100000000001100000000000",--6202
"001101001010000001010000000000000110",--6203
"011100001011000000000000000000000001",--6204
"101110000111111000000001100000000010",--6205
"111110000110010001110001100000000000",--6206
"111110001100011000000010000000000000",--6207
"111110000110001001000001100000000000",--6208
"001011000000000000110000000100101111",--6209
"101001000000000001010000000000000001",--6210
"000101000000000000000001101000011000",--6211
"001101001000000001000000000101101101",--6212
"001101001000000001000000000000000110",--6213
"010000001000000000001111100000000000",--6214
"101001000010000000010000000000000001",--6215
"001100000100000000010010000000000000",--6216
"010011001000000000001111100000000000",--6217
"001101001000000001010000000101101101",--6218
"001111000000000000110000000100010101",--6219
"001101001010000001100000000000000101",--6220
"001111001100000001000000000000000000",--6221
"111110000110010001000001100000000000",--6222
"001111000000000001000000000100010110",--6223
"001111001100000001010000000000000001",--6224
"111110001000010001010010000000000000",--6225
"001111000000000001010000000100010111",--6226
"001111001100000001100000000000000010",--6227
"111110001010010001100010100000000000",--6228
"001101001010000001100000000000000001",--6229
"011111001101000000010000000001010100",--6230
"001111000110000001100000000000000000",--6231
"010010001101000000000000000000011010",--6232
"001101001010000001100000000000000100",--6233
"001101001010000001110000000000000110",--6234
"011010001101000000000000000000000010",--6235
"101001000000000010000000000000000001",--6236
"000101000000000000000001100001011111",--6237
"101000000001111000000100000000000000",--6238
"001111001100000001100000000000000000",--6239
"011100001111000010000000000000000001",--6240
"101110001101111000000011000000000010",--6241
"111110001100010000110011000000000000",--6242
"001111000110000001110000000000000000",--6243
"111110001110011000000011100000000000",--6244
"111110001100001001110011000000000000",--6245
"001111000110000001110000000000000001",--6246
"111110001100001001110011100000000000",--6247
"111110001110000001000011100000000001",--6248
"001111001100000010000000000000000001",--6249
"010110010001000001110000000000001000",--6250
"001111000110000001110000000000000010",--6251
"111110001100001001110011100000000000",--6252
"111110001110000001010011100000000001",--6253
"001111001100000010000000000000000010",--6254
"010110010001000001110000000000000011",--6255
"001011000000000001100000000100101111",--6256
"101001000000000001010000000000000001",--6257
"000101000000000000000001100100111111",--6258
"001111000110000001100000000000000001",--6259
"010010001101000000000000000000011010",--6260
"001101001010000001100000000000000100",--6261
"001101001010000001110000000000000110",--6262
"011010001101000000000000000000000010",--6263
"101001000000000010000000000000000001",--6264
"000101000000000000000001100001111011",--6265
"101000000001111000000100000000000000",--6266
"001111001100000001100000000000000001",--6267
"011100001111000010000000000000000001",--6268
"101110001101111000000011000000000010",--6269
"111110001100010001000011000000000000",--6270
"001111000110000001110000000000000001",--6271
"111110001110011000000011100000000000",--6272
"111110001100001001110011000000000000",--6273
"001111000110000001110000000000000010",--6274
"111110001100001001110011100000000000",--6275
"111110001110000001010011100000000001",--6276
"001111001100000010000000000000000010",--6277
"010110010001000001110000000000001000",--6278
"001111000110000001110000000000000000",--6279
"111110001100001001110011100000000000",--6280
"111110001110000000110011100000000001",--6281
"001111001100000010000000000000000000",--6282
"010110010001000001110000000000000011",--6283
"001011000000000001100000000100101111",--6284
"101001000000000001010000000000000010",--6285
"000101000000000000000001100100111111",--6286
"001111000110000001100000000000000010",--6287
"010010001101000000000000000010101001",--6288
"001101001010000001100000000000000100",--6289
"001101001010000001010000000000000110",--6290
"011010001101000000000000000000000010",--6291
"101001000000000001110000000000000001",--6292
"000101000000000000000001100010010111",--6293
"101000000001111000000011100000000000",--6294
"001111001100000001100000000000000010",--6295
"011100001011000001110000000000000001",--6296
"101110001101111000000011000000000010",--6297
"111110001100010001010010100000000000",--6298
"001111000110000001100000000000000010",--6299
"111110001100011000000011000000000000",--6300
"111110001010001001100010100000000000",--6301
"001111000110000001100000000000000000",--6302
"111110001010001001100011000000000000",--6303
"111110001100000000110001100000000001",--6304
"001111001100000001100000000000000000",--6305
"010110001101000000110000000010010111",--6306
"001111000110000000110000000000000001",--6307
"111110001010001000110001100000000000",--6308
"111110000110000001000001100000000001",--6309
"001111001100000001000000000000000001",--6310
"010110001001000000110000000010010010",--6311
"001011000000000001010000000100101111",--6312
"101001000000000001010000000000000011",--6313
"000101000000000000000001100100111111",--6314
"011111001101000000100000000000011010",--6315
"001101001010000001010000000000000100",--6316
"001111000110000001100000000000000000",--6317
"001111001010000001110000000000000000",--6318
"111110001100001001110011000000000000",--6319
"001111000110000001110000000000000001",--6320
"001111001010000010000000000000000001",--6321
"111110001110001010000011100000000000",--6322
"111110001100000001110011000000000000",--6323
"001111000110000001110000000000000010",--6324
"001111001010000010000000000000000010",--6325
"111110001110001010000011100000000000",--6326
"111110001100000001110011000000000000",--6327
"010110001101000000000000000010000001",--6328
"001111001010000001110000000000000000",--6329
"111110001110001000110001100000000000",--6330
"001111001010000001110000000000000001",--6331
"111110001110001001000010000000000000",--6332
"111110000110000001000001100000000000",--6333
"001111001010000001000000000000000010",--6334
"111110001000001001010010000000000000",--6335
"111110000110000001000001100000000010",--6336
"111110001100011000000010000000000000",--6337
"111110000110001001000001100000000000",--6338
"001011000000000000110000000100101111",--6339
"101001000000000001010000000000000001",--6340
"000101000000000000000001100100111111",--6341
"001111000110000001100000000000000000",--6342
"001111000110000001110000000000000001",--6343
"001111000110000010000000000000000010",--6344
"111110001100001001100100100000000000",--6345
"001101001010000001110000000000000100",--6346
"001111001110000010100000000000000000",--6347
"111110010010001010100100100000000000",--6348
"111110001110001001110101000000000000",--6349
"001111001110000010110000000000000001",--6350
"111110010100001010110101000000000000",--6351
"111110010010000010100100100000000000",--6352
"111110010000001010000101000000000000",--6353
"001111001110000010110000000000000010",--6354
"111110010100001010110101000000000000",--6355
"111110010010000010100100100000000000",--6356
"001101001010000010000000000000000011",--6357
"011100010001000000000000000000000011",--6358
"101110010011111000000011000000000000",--6359
"011110010011000000000000000000001111",--6360
"000101000000000000000001100100111010",--6361
"111110001110001010000101000000000000",--6362
"001101001010000010010000000000001001",--6363
"001111010010000010110000000000000000",--6364
"111110010100001010110101000000000000",--6365
"111110010010000010100100100000000000",--6366
"111110010000001001100100000000000000",--6367
"001111010010000010100000000000000001",--6368
"111110010000001010100100000000000000",--6369
"111110010010000010000100000000000000",--6370
"111110001100001001110011000000000000",--6371
"001111010010000001110000000000000010",--6372
"111110001100001001110011000000000000",--6373
"111110010000000001100011000000000000",--6374
"010010001101000000000000000001010010",--6375
"001111000110000001110000000000000000",--6376
"001111000110000010000000000000000001",--6377
"001111000110000010010000000000000010",--6378
"111110001110001000110101000000000000",--6379
"001111001110000010110000000000000000",--6380
"111110010100001010110101000000000000",--6381
"111110010000001001000101100000000000",--6382
"001111001110000011000000000000000001",--6383
"111110010110001011000101100000000000",--6384
"111110010100000010110101000000000000",--6385
"111110010010001001010101100000000000",--6386
"001111001110000011000000000000000010",--6387
"111110010110001011000101100000000000",--6388
"111110010100000010110101000000000000",--6389
"011100010001000000000000000000000010",--6390
"101110010101111000000011100000000000",--6391
"000101000000000000000001100100001110",--6392
"111110010010001001000101100000000000",--6393
"111110010000001001010110000000000000",--6394
"111110010110000011000101100000000000",--6395
"001101001010000010010000000000001001",--6396
"001111010010000011000000000000000000",--6397
"111110010110001011000101100000000000",--6398
"111110001110001001010110000000000000",--6399
"111110010010001000110100100000000000",--6400
"111110011000000010010100100000000000",--6401
"001111010010000011000000000000000001",--6402
"111110010010001011000100100000000000",--6403
"111110010110000010010100100000000000",--6404
"111110001110001001000011100000000000",--6405
"111110010000001000110100000000000000",--6406
"111110001110000010000011100000000000",--6407
"001111010010000010000000000000000010",--6408
"111110001110001010000011100000000000",--6409
"111110010010000001110011100000000000",--6410
"101111000001110010000011111100000000",--6411
"111110001110001010000011100000000000",--6412
"111110010100000001110011100000000000",--6413
"111110000110001000110100000000000000",--6414
"001111001110000010010000000000000000",--6415
"111110010000001010010100000000000000",--6416
"111110001000001001000100100000000000",--6417
"001111001110000010100000000000000001",--6418
"111110010010001010100100100000000000",--6419
"111110010000000010010100000000000000",--6420
"111110001010001001010100100000000000",--6421
"001111001110000010100000000000000010",--6422
"111110010010001010100100100000000000",--6423
"111110010000000010010100000000000000",--6424
"011100010001000000000000000000000011",--6425
"101110010001111000000001100000000000",--6426
"011111001101000000110000000000010000",--6427
"000101000000000000000001100100101011",--6428
"111110001000001001010100100000000000",--6429
"001101001010000001110000000000001001",--6430
"001111001110000010100000000000000000",--6431
"111110010010001010100100100000000000",--6432
"111110010000000010010100000000000000",--6433
"111110001010001000110010100000000000",--6434
"001111001110000010010000000000000001",--6435
"111110001010001010010010100000000000",--6436
"111110010000000001010010100000000000",--6437
"111110000110001001000001100000000000",--6438
"001111001110000001000000000000000010",--6439
"111110000110001001000001100000000000",--6440
"111110001010000000110001100000000000",--6441
"011111001101000000110000000000000001",--6442
"111110000110010000010001100000000000",--6443
"111110001110001001110010000000000000",--6444
"111110001100001000110001100000000000",--6445
"111110001000010000110001100000000000",--6446
"010110000111000000000000000000001010",--6447
"111110000110100000000001100000000000",--6448
"001101001010000001010000000000000110",--6449
"011100001011000000000000000000000001",--6450
"101110000111111000000001100000000010",--6451
"111110000110010001110001100000000000",--6452
"111110001100011000000010000000000000",--6453
"111110000110001001000001100000000000",--6454
"001011000000000000110000000100101111",--6455
"101001000000000001010000000000000001",--6456
"000101000000000000000001100100111111",--6457
"001101001000000001000000000101101101",--6458
"001101001000000001000000000000000110",--6459
"010000001000000000001111100000000000",--6460
"101001000010000000010000000000000001",--6461
"000101000000000000000001011101010010",--6462
"001111000000000000110000000100101111",--6463
"001001111100000000110000000000000000",--6464
"001001111100000000101111111111111111",--6465
"001001111100000000011111111111111110",--6466
"010110000111000000000000000011001111",--6467
"001111000000000001000000000100101101",--6468
"010110001001000000110000000011001101",--6469
"101111001001110001000011110000100011",--6470
"101111001001100001001101011100001010",--6471
"111110000110000001000001100000000000",--6472
"001111000110000001000000000000000000",--6473
"111110001000001000110010000000000000",--6474
"001111000000000001010000000100010101",--6475
"111110001000000001010010000000000000",--6476
"001111000110000001010000000000000001",--6477
"111110001010001000110010100000000000",--6478
"001111000000000001100000000100010110",--6479
"111110001010000001100010100000000000",--6480
"001111000110000001100000000000000010",--6481
"111110001100001000110011000000000000",--6482
"001111000000000001110000000100010111",--6483
"111110001100000001110011000000000000",--6484
"001101000100000001100000000000000000",--6485
"001001111100000001011111111111111101",--6486
"001001111100000001001111111111111100",--6487
"001011111100000001101111111111111011",--6488
"001011111100000001011111111111111010",--6489
"001011111100000001001111111111111001",--6490
"001011111100000000111111111111111000",--6491
"010011001101000000000000000010101010",--6492
"001101001100000001100000000101101101",--6493
"001101001100000001110000000000000101",--6494
"001111001110000001110000000000000000",--6495
"111110001000010001110011100000000000",--6496
"001111001110000010000000000000000001",--6497
"111110001010010010000100000000000000",--6498
"001111001110000010010000000000000010",--6499
"111110001100010010010100100000000000",--6500
"001101001100000001110000000000000001",--6501
"011111001111000000010000000000010000",--6502
"101110001111111000000011100000000001",--6503
"001101001100000001110000000000000100",--6504
"001111001110000010100000000000000000",--6505
"010110010101000001110000000000001001",--6506
"101110010001111000000011100000000001",--6507
"001111001110000010000000000000000001",--6508
"010110010001000001110000000000000110",--6509
"101110010011111000000011100000000001",--6510
"001111001110000010000000000000000010",--6511
"010110010001000001110000000000000011",--6512
"001101001100000001100000000000000110",--6513
"011100001101000000000000000010100000",--6514
"000101000000000000000001100110101100",--6515
"001101001100000001100000000000000110",--6516
"011100001101000000000000000000110110",--6517
"000101000000000000000001101000010011",--6518
"011111001111000000100000000000001111",--6519
"001101001100000001110000000000000100",--6520
"001111001110000010100000000000000000",--6521
"111110010100001001110011100000000000",--6522
"001111001110000010100000000000000001",--6523
"111110010100001010000100000000000000",--6524
"111110001110000010000011100000000000",--6525
"001111001110000010000000000000000010",--6526
"111110010000001010010100000000000000",--6527
"111110001110000010000011100000000000",--6528
"001101001100000001100000000000000110",--6529
"011010001111000000000000000000000010",--6530
"011111001101000000010000000000101000",--6531
"000101000000000000000001101000010011",--6532
"011100001101000000000000000000100110",--6533
"000101000000000000000001101000010011",--6534
"111110001110001001110101000000000000",--6535
"001101001100000010000000000000000100",--6536
"001111010000000010110000000000000000",--6537
"111110010100001010110101000000000000",--6538
"111110010000001010000101100000000000",--6539
"001111010000000011000000000000000001",--6540
"111110010110001011000101100000000000",--6541
"111110010100000010110101000000000000",--6542
"111110010010001010010101100000000000",--6543
"001111010000000011000000000000000010",--6544
"111110010110001011000101100000000000",--6545
"111110010100000010110101000000000000",--6546
"001101001100000010000000000000000011",--6547
"011100010001000000000000000000000011",--6548
"101110010101111000000011100000000000",--6549
"011111001111000000110000000000010000",--6550
"000101000000000000000001100110100110",--6551
"111110010000001010010101100000000000",--6552
"001101001100000010000000000000001001",--6553
"001111010000000011000000000000000000",--6554
"111110010110001011000101100000000000",--6555
"111110010100000010110101000000000000",--6556
"111110010010001001110100100000000000",--6557
"001111010000000010110000000000000001",--6558
"111110010010001010110100100000000000",--6559
"111110010100000010010100100000000000",--6560
"111110001110001010000011100000000000",--6561
"001111010000000010000000000000000010",--6562
"111110001110001010000011100000000000",--6563
"111110010010000001110011100000000000",--6564
"011111001111000000110000000000000001",--6565
"111110001110010000010011100000000000",--6566
"001101001100000001100000000000000110",--6567
"011010001111000000000000000000000010",--6568
"011111001101000000010000000000000010",--6569
"000101000000000000000001101000010011",--6570
"010000001101000000000000000001100111",--6571
"001101000100000001100000000000000001",--6572
"010011001101000000000000000001011001",--6573
"001101001100000001100000000101101101",--6574
"001101001100000001110000000000000101",--6575
"001111001110000001110000000000000000",--6576
"111110001000010001110011100000000000",--6577
"001111001110000010000000000000000001",--6578
"111110001010010010000100000000000000",--6579
"001111001110000010010000000000000010",--6580
"111110001100010010010100100000000000",--6581
"001101001100000001110000000000000001",--6582
"011111001111000000010000000000010000",--6583
"101110001111111000000011100000000001",--6584
"001101001100000001110000000000000100",--6585
"001111001110000010100000000000000000",--6586
"010110010101000001110000000000001001",--6587
"101110010001111000000011100000000001",--6588
"001111001110000010000000000000000001",--6589
"010110010001000001110000000000000110",--6590
"101110010011111000000011100000000001",--6591
"001111001110000010000000000000000010",--6592
"010110010001000001110000000000000011",--6593
"001101001100000001100000000000000110",--6594
"011100001101000000000000000001001111",--6595
"000101000000000000000001100111111101",--6596
"001101001100000001100000000000000110",--6597
"011100001101000000000000000000110110",--6598
"000101000000000000000001101000010011",--6599
"011111001111000000100000000000001111",--6600
"001101001100000001110000000000000100",--6601
"001111001110000010100000000000000000",--6602
"111110010100001001110011100000000000",--6603
"001111001110000010100000000000000001",--6604
"111110010100001010000100000000000000",--6605
"111110001110000010000011100000000000",--6606
"001111001110000010000000000000000010",--6607
"111110010000001010010100000000000000",--6608
"111110001110000010000011100000000000",--6609
"001101001100000001100000000000000110",--6610
"011010001111000000000000000000000010",--6611
"011111001101000000010000000000101000",--6612
"000101000000000000000001101000010011",--6613
"011100001101000000000000000000100110",--6614
"000101000000000000000001101000010011",--6615
"111110001110001001110101000000000000",--6616
"001101001100000010000000000000000100",--6617
"001111010000000010110000000000000000",--6618
"111110010100001010110101000000000000",--6619
"111110010000001010000101100000000000",--6620
"001111010000000011000000000000000001",--6621
"111110010110001011000101100000000000",--6622
"111110010100000010110101000000000000",--6623
"111110010010001010010101100000000000",--6624
"001111010000000011000000000000000010",--6625
"111110010110001011000101100000000000",--6626
"111110010100000010110101000000000000",--6627
"001101001100000010000000000000000011",--6628
"011100010001000000000000000000000011",--6629
"101110010101111000000011100000000000",--6630
"011111001111000000110000000000010000",--6631
"000101000000000000000001100111110111",--6632
"111110010000001010010101100000000000",--6633
"001101001100000010000000000000001001",--6634
"001111010000000011000000000000000000",--6635
"111110010110001011000101100000000000",--6636
"111110010100000010110101000000000000",--6637
"111110010010001001110100100000000000",--6638
"001111010000000010110000000000000001",--6639
"111110010010001010110100100000000000",--6640
"111110010100000010010100100000000000",--6641
"111110001110001010000011100000000000",--6642
"001111010000000010000000000000000010",--6643
"111110001110001010000011100000000000",--6644
"111110010010000001110011100000000000",--6645
"011111001111000000110000000000000001",--6646
"111110001110010000010011100000000000",--6647
"001101001100000001100000000000000110",--6648
"011010001111000000000000000000000010",--6649
"011111001101000000010000000000000010",--6650
"000101000000000000000001101000010011",--6651
"010000001101000000000000000000010110",--6652
"101001000000000000010000000000000010",--6653
"101110001001111000000001100000000000",--6654
"101110001011111000000010000000000000",--6655
"101110001101111000000010100000000000",--6656
"001001111100000111111111111111110111",--6657
"101001111100010111100000000000001010",--6658
"000111000000000000000000011110001000",--6659
"101001111100000111100000000000001010",--6660
"001101111100000111111111111111110111",--6661
"010000000011000000000000000000001100",--6662
"001111111100000000111111111111111000",--6663
"001011000000000000110000000100101101",--6664
"001111111100000000111111111111111001",--6665
"001011000000000000110000000100101010",--6666
"001111111100000000111111111111111010",--6667
"001011000000000000110000000100101011",--6668
"001111111100000000111111111111111011",--6669
"001011000000000000110000000100101100",--6670
"001101111100000000011111111111111100",--6671
"001001000000000000010000000100101001",--6672
"001101111100000000011111111111111101",--6673
"001001000000000000010000000100101110",--6674
"001101111100000000011111111111111110",--6675
"101001000010000000010000000000000001",--6676
"001101111100000000101111111111111111",--6677
"001101111100000000110000000000000000",--6678
"000101000000000000000001011101010010",--6679
"001111000000000000110000000100101111",--6680
"001001111100000000110000000000000000",--6681
"001001111100000000101111111111111111",--6682
"001001111100000000011111111111111110",--6683
"010110000111000000000000000100100000",--6684
"001111000000000001000000000100101101",--6685
"010110001001000000110000000100011110",--6686
"101111001001110001000011110000100011",--6687
"101111001001100001001101011100001010",--6688
"111110000110000001000001100000000000",--6689
"001111000110000001000000000000000000",--6690
"111110001000001000110010000000000000",--6691
"001111000000000001010000000100010101",--6692
"111110001000000001010010000000000000",--6693
"001111000110000001010000000000000001",--6694
"111110001010001000110010100000000000",--6695
"001111000000000001100000000100010110",--6696
"111110001010000001100010100000000000",--6697
"001111000110000001100000000000000010",--6698
"111110001100001000110011000000000000",--6699
"001111000000000001110000000100010111",--6700
"111110001100000001110011000000000000",--6701
"001101000100000001100000000000000000",--6702
"001001111100000001011111111111111101",--6703
"001001111100000001001111111111111100",--6704
"001011111100000001101111111111111011",--6705
"001011111100000001011111111111111010",--6706
"001011111100000001001111111111111001",--6707
"001011111100000000111111111111111000",--6708
"010011001101000000000000000011111011",--6709
"001101001100000001100000000101101101",--6710
"001101001100000001110000000000000101",--6711
"001111001110000001110000000000000000",--6712
"111110001000010001110011100000000000",--6713
"001111001110000010000000000000000001",--6714
"111110001010010010000100000000000000",--6715
"001111001110000010010000000000000010",--6716
"111110001100010010010100100000000000",--6717
"001101001100000001110000000000000001",--6718
"011111001111000000010000000000010000",--6719
"101110001111111000000011100000000001",--6720
"001101001100000001110000000000000100",--6721
"001111001110000010100000000000000000",--6722
"010110010101000001110000000000001001",--6723
"101110010001111000000011100000000001",--6724
"001111001110000010000000000000000001",--6725
"010110010001000001110000000000000110",--6726
"101110010011111000000011100000000001",--6727
"001111001110000010000000000000000010",--6728
"010110010001000001110000000000000011",--6729
"001101001100000001100000000000000110",--6730
"011100001101000000000000000011110001",--6731
"000101000000000000000001101010000101",--6732
"001101001100000001100000000000000110",--6733
"011100001101000000000000000000110110",--6734
"000101000000000000000001101100111101",--6735
"011111001111000000100000000000001111",--6736
"001101001100000001110000000000000100",--6737
"001111001110000010100000000000000000",--6738
"111110010100001001110011100000000000",--6739
"001111001110000010100000000000000001",--6740
"111110010100001010000100000000000000",--6741
"111110001110000010000011100000000000",--6742
"001111001110000010000000000000000010",--6743
"111110010000001010010100000000000000",--6744
"111110001110000010000011100000000000",--6745
"001101001100000001100000000000000110",--6746
"011010001111000000000000000000000010",--6747
"011111001101000000010000000000101000",--6748
"000101000000000000000001101100111101",--6749
"011100001101000000000000000000100110",--6750
"000101000000000000000001101100111101",--6751
"111110001110001001110101000000000000",--6752
"001101001100000010000000000000000100",--6753
"001111010000000010110000000000000000",--6754
"111110010100001010110101000000000000",--6755
"111110010000001010000101100000000000",--6756
"001111010000000011000000000000000001",--6757
"111110010110001011000101100000000000",--6758
"111110010100000010110101000000000000",--6759
"111110010010001010010101100000000000",--6760
"001111010000000011000000000000000010",--6761
"111110010110001011000101100000000000",--6762
"111110010100000010110101000000000000",--6763
"001101001100000010000000000000000011",--6764
"011100010001000000000000000000000011",--6765
"101110010101111000000011100000000000",--6766
"011111001111000000110000000000010000",--6767
"000101000000000000000001101001111111",--6768
"111110010000001010010101100000000000",--6769
"001101001100000010000000000000001001",--6770
"001111010000000011000000000000000000",--6771
"111110010110001011000101100000000000",--6772
"111110010100000010110101000000000000",--6773
"111110010010001001110100100000000000",--6774
"001111010000000010110000000000000001",--6775
"111110010010001010110100100000000000",--6776
"111110010100000010010100100000000000",--6777
"111110001110001010000011100000000000",--6778
"001111010000000010000000000000000010",--6779
"111110001110001010000011100000000000",--6780
"111110010010000001110011100000000000",--6781
"011111001111000000110000000000000001",--6782
"111110001110010000010011100000000000",--6783
"001101001100000001100000000000000110",--6784
"011010001111000000000000000000000010",--6785
"011111001101000000010000000000000010",--6786
"000101000000000000000001101100111101",--6787
"010000001101000000000000000010111000",--6788
"001101000100000001100000000000000001",--6789
"010011001101000000000000000010101010",--6790
"001101001100000001100000000101101101",--6791
"001101001100000001110000000000000101",--6792
"001111001110000001110000000000000000",--6793
"111110001000010001110011100000000000",--6794
"001111001110000010000000000000000001",--6795
"111110001010010010000100000000000000",--6796
"001111001110000010010000000000000010",--6797
"111110001100010010010100100000000000",--6798
"001101001100000001110000000000000001",--6799
"011111001111000000010000000000010000",--6800
"101110001111111000000011100000000001",--6801
"001101001100000001110000000000000100",--6802
"001111001110000010100000000000000000",--6803
"010110010101000001110000000000001001",--6804
"101110010001111000000011100000000001",--6805
"001111001110000010000000000000000001",--6806
"010110010001000001110000000000000110",--6807
"101110010011111000000011100000000001",--6808
"001111001110000010000000000000000010",--6809
"010110010001000001110000000000000011",--6810
"001101001100000001100000000000000110",--6811
"011100001101000000000000000010100000",--6812
"000101000000000000000001101011010110",--6813
"001101001100000001100000000000000110",--6814
"011100001101000000000000000000110110",--6815
"000101000000000000000001101100111101",--6816
"011111001111000000100000000000001111",--6817
"001101001100000001110000000000000100",--6818
"001111001110000010100000000000000000",--6819
"111110010100001001110011100000000000",--6820
"001111001110000010100000000000000001",--6821
"111110010100001010000100000000000000",--6822
"111110001110000010000011100000000000",--6823
"001111001110000010000000000000000010",--6824
"111110010000001010010100000000000000",--6825
"111110001110000010000011100000000000",--6826
"001101001100000001100000000000000110",--6827
"011010001111000000000000000000000010",--6828
"011111001101000000010000000000101000",--6829
"000101000000000000000001101100111101",--6830
"011100001101000000000000000000100110",--6831
"000101000000000000000001101100111101",--6832
"111110001110001001110101000000000000",--6833
"001101001100000010000000000000000100",--6834
"001111010000000010110000000000000000",--6835
"111110010100001010110101000000000000",--6836
"111110010000001010000101100000000000",--6837
"001111010000000011000000000000000001",--6838
"111110010110001011000101100000000000",--6839
"111110010100000010110101000000000000",--6840
"111110010010001010010101100000000000",--6841
"001111010000000011000000000000000010",--6842
"111110010110001011000101100000000000",--6843
"111110010100000010110101000000000000",--6844
"001101001100000010000000000000000011",--6845
"011100010001000000000000000000000011",--6846
"101110010101111000000011100000000000",--6847
"011111001111000000110000000000010000",--6848
"000101000000000000000001101011010000",--6849
"111110010000001010010101100000000000",--6850
"001101001100000010000000000000001001",--6851
"001111010000000011000000000000000000",--6852
"111110010110001011000101100000000000",--6853
"111110010100000010110101000000000000",--6854
"111110010010001001110100100000000000",--6855
"001111010000000010110000000000000001",--6856
"111110010010001010110100100000000000",--6857
"111110010100000010010100100000000000",--6858
"111110001110001010000011100000000000",--6859
"001111010000000010000000000000000010",--6860
"111110001110001010000011100000000000",--6861
"111110010010000001110011100000000000",--6862
"011111001111000000110000000000000001",--6863
"111110001110010000010011100000000000",--6864
"001101001100000001100000000000000110",--6865
"011010001111000000000000000000000010",--6866
"011111001101000000010000000000000010",--6867
"000101000000000000000001101100111101",--6868
"010000001101000000000000000001100111",--6869
"001101000100000001100000000000000010",--6870
"010011001101000000000000000001011001",--6871
"001101001100000001100000000101101101",--6872
"001101001100000001110000000000000101",--6873
"001111001110000001110000000000000000",--6874
"111110001000010001110011100000000000",--6875
"001111001110000010000000000000000001",--6876
"111110001010010010000100000000000000",--6877
"001111001110000010010000000000000010",--6878
"111110001100010010010100100000000000",--6879
"001101001100000001110000000000000001",--6880
"011111001111000000010000000000010000",--6881
"101110001111111000000011100000000001",--6882
"001101001100000001110000000000000100",--6883
"001111001110000010100000000000000000",--6884
"010110010101000001110000000000001001",--6885
"101110010001111000000011100000000001",--6886
"001111001110000010000000000000000001",--6887
"010110010001000001110000000000000110",--6888
"101110010011111000000011100000000001",--6889
"001111001110000010000000000000000010",--6890
"010110010001000001110000000000000011",--6891
"001101001100000001100000000000000110",--6892
"011100001101000000000000000001001111",--6893
"000101000000000000000001101100100111",--6894
"001101001100000001100000000000000110",--6895
"011100001101000000000000000000110110",--6896
"000101000000000000000001101100111101",--6897
"011111001111000000100000000000001111",--6898
"001101001100000001110000000000000100",--6899
"001111001110000010100000000000000000",--6900
"111110010100001001110011100000000000",--6901
"001111001110000010100000000000000001",--6902
"111110010100001010000100000000000000",--6903
"111110001110000010000011100000000000",--6904
"001111001110000010000000000000000010",--6905
"111110010000001010010100000000000000",--6906
"111110001110000010000011100000000000",--6907
"001101001100000001100000000000000110",--6908
"011010001111000000000000000000000010",--6909
"011111001101000000010000000000101000",--6910
"000101000000000000000001101100111101",--6911
"011100001101000000000000000000100110",--6912
"000101000000000000000001101100111101",--6913
"111110001110001001110101000000000000",--6914
"001101001100000010000000000000000100",--6915
"001111010000000010110000000000000000",--6916
"111110010100001010110101000000000000",--6917
"111110010000001010000101100000000000",--6918
"001111010000000011000000000000000001",--6919
"111110010110001011000101100000000000",--6920
"111110010100000010110101000000000000",--6921
"111110010010001010010101100000000000",--6922
"001111010000000011000000000000000010",--6923
"111110010110001011000101100000000000",--6924
"111110010100000010110101000000000000",--6925
"001101001100000010000000000000000011",--6926
"011100010001000000000000000000000011",--6927
"101110010101111000000011100000000000",--6928
"011111001111000000110000000000010000",--6929
"000101000000000000000001101100100001",--6930
"111110010000001010010101100000000000",--6931
"001101001100000010000000000000001001",--6932
"001111010000000011000000000000000000",--6933
"111110010110001011000101100000000000",--6934
"111110010100000010110101000000000000",--6935
"111110010010001001110100100000000000",--6936
"001111010000000010110000000000000001",--6937
"111110010010001010110100100000000000",--6938
"111110010100000010010100100000000000",--6939
"111110001110001010000011100000000000",--6940
"001111010000000010000000000000000010",--6941
"111110001110001010000011100000000000",--6942
"111110010010000001110011100000000000",--6943
"011111001111000000110000000000000001",--6944
"111110001110010000010011100000000000",--6945
"001101001100000001100000000000000110",--6946
"011010001111000000000000000000000010",--6947
"011111001101000000010000000000000010",--6948
"000101000000000000000001101100111101",--6949
"010000001101000000000000000000010110",--6950
"101001000000000000010000000000000011",--6951
"101110001001111000000001100000000000",--6952
"101110001011111000000010000000000000",--6953
"101110001101111000000010100000000000",--6954
"001001111100000111111111111111110111",--6955
"101001111100010111100000000000001010",--6956
"000111000000000000000000011110001000",--6957
"101001111100000111100000000000001010",--6958
"001101111100000111111111111111110111",--6959
"010000000011000000000000000000001100",--6960
"001111111100000000111111111111111000",--6961
"001011000000000000110000000100101101",--6962
"001111111100000000111111111111111001",--6963
"001011000000000000110000000100101010",--6964
"001111111100000000111111111111111010",--6965
"001011000000000000110000000100101011",--6966
"001111111100000000111111111111111011",--6967
"001011000000000000110000000100101100",--6968
"001101111100000000011111111111111100",--6969
"001001000000000000010000000100101001",--6970
"001101111100000000011111111111111101",--6971
"001001000000000000010000000100101110",--6972
"001101111100000000011111111111111110",--6973
"101001000010000000010000000000000001",--6974
"001101111100000000111111111111111111",--6975
"001100000110000000010001000000000000",--6976
"010011000100000000001111100000000000",--6977
"001101000100000001000000000101101101",--6978
"001111000000000000110000000100010101",--6979
"001101001000000001010000000000000101",--6980
"001111001010000001000000000000000000",--6981
"111110000110010001000001100000000000",--6982
"001111000000000001000000000100010110",--6983
"001111001010000001010000000000000001",--6984
"111110001000010001010010000000000000",--6985
"001111000000000001010000000100010111",--6986
"001111001010000001100000000000000010",--6987
"111110001010010001100010100000000000",--6988
"001101001000000001010000000000000001",--6989
"011111001011000000010000000001010101",--6990
"001101111100000001010000000000000000",--6991
"001111001010000001100000000000000000",--6992
"010010001101000000000000000000011010",--6993
"001101001000000001100000000000000100",--6994
"001101001000000001110000000000000110",--6995
"011010001101000000000000000000000010",--6996
"101001000000000010000000000000000001",--6997
"000101000000000000000001101101011000",--6998
"101000000001111000000100000000000000",--6999
"001111001100000001100000000000000000",--7000
"011100001111000010000000000000000001",--7001
"101110001101111000000011000000000010",--7002
"111110001100010000110011000000000000",--7003
"001111001010000001110000000000000000",--7004
"111110001110011000000011100000000000",--7005
"111110001100001001110011000000000000",--7006
"001111001010000001110000000000000001",--7007
"111110001100001001110011100000000000",--7008
"111110001110000001000011100000000001",--7009
"001111001100000010000000000000000001",--7010
"010110010001000001110000000000001000",--7011
"001111001010000001110000000000000010",--7012
"111110001100001001110011100000000000",--7013
"111110001110000001010011100000000001",--7014
"001111001100000010000000000000000010",--7015
"010110010001000001110000000000000011",--7016
"001011000000000001100000000100101111",--7017
"101001000000000001000000000000000001",--7018
"000101000000000000000001110000111110",--7019
"001111001010000001100000000000000001",--7020
"010010001101000000000000000000011010",--7021
"001101001000000001100000000000000100",--7022
"001101001000000001110000000000000110",--7023
"011010001101000000000000000000000010",--7024
"101001000000000010000000000000000001",--7025
"000101000000000000000001101101110100",--7026
"101000000001111000000100000000000000",--7027
"001111001100000001100000000000000001",--7028
"011100001111000010000000000000000001",--7029
"101110001101111000000011000000000010",--7030
"111110001100010001000011000000000000",--7031
"001111001010000001110000000000000001",--7032
"111110001110011000000011100000000000",--7033
"111110001100001001110011000000000000",--7034
"001111001010000001110000000000000010",--7035
"111110001100001001110011100000000000",--7036
"111110001110000001010011100000000001",--7037
"001111001100000010000000000000000010",--7038
"010110010001000001110000000000001000",--7039
"001111001010000001110000000000000000",--7040
"111110001100001001110011100000000000",--7041
"111110001110000000110011100000000001",--7042
"001111001100000010000000000000000000",--7043
"010110010001000001110000000000000011",--7044
"001011000000000001100000000100101111",--7045
"101001000000000001000000000000000010",--7046
"000101000000000000000001110000111110",--7047
"001111001010000001100000000000000010",--7048
"010010001101000000000000000010101011",--7049
"001101001000000001100000000000000100",--7050
"001101001000000001000000000000000110",--7051
"011010001101000000000000000000000010",--7052
"101001000000000001110000000000000001",--7053
"000101000000000000000001101110010000",--7054
"101000000001111000000011100000000000",--7055
"001111001100000001100000000000000010",--7056
"011100001001000001110000000000000001",--7057
"101110001101111000000011000000000010",--7058
"111110001100010001010010100000000000",--7059
"001111001010000001100000000000000010",--7060
"111110001100011000000011000000000000",--7061
"111110001010001001100010100000000000",--7062
"001111001010000001100000000000000000",--7063
"111110001010001001100011000000000000",--7064
"111110001100000000110001100000000001",--7065
"001111001100000001100000000000000000",--7066
"010110001101000000110000000010011001",--7067
"001111001010000000110000000000000001",--7068
"111110001010001000110001100000000000",--7069
"111110000110000001000001100000000001",--7070
"001111001100000001000000000000000001",--7071
"010110001001000000110000000010010100",--7072
"001011000000000001010000000100101111",--7073
"101001000000000001000000000000000011",--7074
"000101000000000000000001110000111110",--7075
"011111001011000000100000000000011011",--7076
"001101001000000001000000000000000100",--7077
"001101111100000001010000000000000000",--7078
"001111001010000001100000000000000000",--7079
"001111001000000001110000000000000000",--7080
"111110001100001001110011000000000000",--7081
"001111001010000001110000000000000001",--7082
"001111001000000010000000000000000001",--7083
"111110001110001010000011100000000000",--7084
"111110001100000001110011000000000000",--7085
"001111001010000001110000000000000010",--7086
"001111001000000010000000000000000010",--7087
"111110001110001010000011100000000000",--7088
"111110001100000001110011000000000000",--7089
"010110001101000000000000000010000010",--7090
"001111001000000001110000000000000000",--7091
"111110001110001000110001100000000000",--7092
"001111001000000001110000000000000001",--7093
"111110001110001001000010000000000000",--7094
"111110000110000001000001100000000000",--7095
"001111001000000001000000000000000010",--7096
"111110001000001001010010000000000000",--7097
"111110000110000001000001100000000010",--7098
"111110001100011000000010000000000000",--7099
"111110000110001001000001100000000000",--7100
"001011000000000000110000000100101111",--7101
"101001000000000001000000000000000001",--7102
"000101000000000000000001110000111110",--7103
"001101111100000001100000000000000000",--7104
"001111001100000001100000000000000000",--7105
"001111001100000001110000000000000001",--7106
"001111001100000010000000000000000010",--7107
"111110001100001001100100100000000000",--7108
"001101001000000001110000000000000100",--7109
"001111001110000010100000000000000000",--7110
"111110010010001010100100100000000000",--7111
"111110001110001001110101000000000000",--7112
"001111001110000010110000000000000001",--7113
"111110010100001010110101000000000000",--7114
"111110010010000010100100100000000000",--7115
"111110010000001010000101000000000000",--7116
"001111001110000010110000000000000010",--7117
"111110010100001010110101000000000000",--7118
"111110010010000010100100100000000000",--7119
"001101001000000010000000000000000011",--7120
"011100010001000000000000000000000011",--7121
"101110010011111000000011000000000000",--7122
"011110010011000000000000000000001111",--7123
"000101000000000000000001110000110101",--7124
"111110001110001010000101000000000000",--7125
"001101001000000010010000000000001001",--7126
"001111010010000010110000000000000000",--7127
"111110010100001010110101000000000000",--7128
"111110010010000010100100100000000000",--7129
"111110010000001001100100000000000000",--7130
"001111010010000010100000000000000001",--7131
"111110010000001010100100000000000000",--7132
"111110010010000010000100000000000000",--7133
"111110001100001001110011000000000000",--7134
"001111010010000001110000000000000010",--7135
"111110001100001001110011000000000000",--7136
"111110010000000001100011000000000000",--7137
"010010001101000000000000000001010010",--7138
"001111001100000001110000000000000000",--7139
"001111001100000010000000000000000001",--7140
"001111001100000010010000000000000010",--7141
"111110001110001000110101000000000000",--7142
"001111001110000010110000000000000000",--7143
"111110010100001010110101000000000000",--7144
"111110010000001001000101100000000000",--7145
"001111001110000011000000000000000001",--7146
"111110010110001011000101100000000000",--7147
"111110010100000010110101000000000000",--7148
"111110010010001001010101100000000000",--7149
"001111001110000011000000000000000010",--7150
"111110010110001011000101100000000000",--7151
"111110010100000010110101000000000000",--7152
"011100010001000000000000000000000010",--7153
"101110010101111000000011100000000000",--7154
"000101000000000000000001110000001001",--7155
"111110010010001001000101100000000000",--7156
"111110010000001001010110000000000000",--7157
"111110010110000011000101100000000000",--7158
"001101001000000010010000000000001001",--7159
"001111010010000011000000000000000000",--7160
"111110010110001011000101100000000000",--7161
"111110001110001001010110000000000000",--7162
"111110010010001000110100100000000000",--7163
"111110011000000010010100100000000000",--7164
"001111010010000011000000000000000001",--7165
"111110010010001011000100100000000000",--7166
"111110010110000010010100100000000000",--7167
"111110001110001001000011100000000000",--7168
"111110010000001000110100000000000000",--7169
"111110001110000010000011100000000000",--7170
"001111010010000010000000000000000010",--7171
"111110001110001010000011100000000000",--7172
"111110010010000001110011100000000000",--7173
"101111000001110010000011111100000000",--7174
"111110001110001010000011100000000000",--7175
"111110010100000001110011100000000000",--7176
"111110000110001000110100000000000000",--7177
"001111001110000010010000000000000000",--7178
"111110010000001010010100000000000000",--7179
"111110001000001001000100100000000000",--7180
"001111001110000010100000000000000001",--7181
"111110010010001010100100100000000000",--7182
"111110010000000010010100000000000000",--7183
"111110001010001001010100100000000000",--7184
"001111001110000010100000000000000010",--7185
"111110010010001010100100100000000000",--7186
"111110010000000010010100000000000000",--7187
"011100010001000000000000000000000011",--7188
"101110010001111000000001100000000000",--7189
"011111001011000000110000000000010000",--7190
"000101000000000000000001110000100110",--7191
"111110001000001001010100100000000000",--7192
"001101001000000001110000000000001001",--7193
"001111001110000010100000000000000000",--7194
"111110010010001010100100100000000000",--7195
"111110010000000010010100000000000000",--7196
"111110001010001000110010100000000000",--7197
"001111001110000010010000000000000001",--7198
"111110001010001010010010100000000000",--7199
"111110010000000001010010100000000000",--7200
"111110000110001001000001100000000000",--7201
"001111001110000001000000000000000010",--7202
"111110000110001001000001100000000000",--7203
"111110001010000000110001100000000000",--7204
"011111001011000000110000000000000001",--7205
"111110000110010000010001100000000000",--7206
"111110001110001001110010000000000000",--7207
"111110001100001000110001100000000000",--7208
"111110001000010000110001100000000000",--7209
"010110000111000000000000000000001010",--7210
"111110000110100000000001100000000000",--7211
"001101001000000001000000000000000110",--7212
"011100001001000000000000000000000001",--7213
"101110000111111000000001100000000010",--7214
"111110000110010001110001100000000000",--7215
"111110001100011000000010000000000000",--7216
"111110000110001001000001100000000000",--7217
"001011000000000000110000000100101111",--7218
"101001000000000001000000000000000001",--7219
"000101000000000000000001110000111110",--7220
"001101000100000000100000000101101101",--7221
"001101000100000000100000000000000110",--7222
"010000000100000000001111100000000000",--7223
"101001000010000000010000000000000001",--7224
"001101111100000000100000000000000000",--7225
"101000000111111000001101100000000000",--7226
"101000000101111000000001100000000000",--7227
"101000110111111000000001000000000000",--7228
"000101000000000000000001011101010010",--7229
"001111000000000000110000000100101111",--7230
"001001111100000000011111111111111101",--7231
"010110000111000000000000000011010001",--7232
"001111000000000001000000000100101101",--7233
"010110001001000000110000000011001111",--7234
"101111001001110001000011110000100011",--7235
"101111001001100001001101011100001010",--7236
"111110000110000001000001100000000000",--7237
"001101111100000001010000000000000000",--7238
"001111001010000001000000000000000000",--7239
"111110001000001000110010000000000000",--7240
"001111000000000001010000000100010101",--7241
"111110001000000001010010000000000000",--7242
"001111001010000001010000000000000001",--7243
"111110001010001000110010100000000000",--7244
"001111000000000001100000000100010110",--7245
"111110001010000001100010100000000000",--7246
"001111001010000001100000000000000010",--7247
"111110001100001000110011000000000000",--7248
"001111000000000001110000000100010111",--7249
"111110001100000001110011000000000000",--7250
"001101000110000001100000000000000000",--7251
"001001111100000001001111111111111100",--7252
"001001111100000000101111111111111011",--7253
"001011111100000001101111111111111010",--7254
"001011111100000001011111111111111001",--7255
"001011111100000001001111111111111000",--7256
"001011111100000000111111111111110111",--7257
"010011001101000000000000000010101011",--7258
"001101001100000001100000000101101101",--7259
"001101001100000001110000000000000101",--7260
"001111001110000001110000000000000000",--7261
"111110001000010001110011100000000000",--7262
"001111001110000010000000000000000001",--7263
"111110001010010010000100000000000000",--7264
"001111001110000010010000000000000010",--7265
"111110001100010010010100100000000000",--7266
"001101001100000001110000000000000001",--7267
"011111001111000000010000000000010000",--7268
"101110001111111000000011100000000001",--7269
"001101001100000001110000000000000100",--7270
"001111001110000010100000000000000000",--7271
"010110010101000001110000000000001001",--7272
"101110010001111000000011100000000001",--7273
"001111001110000010000000000000000001",--7274
"010110010001000001110000000000000110",--7275
"101110010011111000000011100000000001",--7276
"001111001110000010000000000000000010",--7277
"010110010001000001110000000000000011",--7278
"001101001100000001100000000000000110",--7279
"011100001101000000000000000010100001",--7280
"000101000000000000000001110010101010",--7281
"001101001100000001100000000000000110",--7282
"011100001101000000000000000000110110",--7283
"000101000000000000000001110100010010",--7284
"011111001111000000100000000000001111",--7285
"001101001100000001110000000000000100",--7286
"001111001110000010100000000000000000",--7287
"111110010100001001110011100000000000",--7288
"001111001110000010100000000000000001",--7289
"111110010100001010000100000000000000",--7290
"111110001110000010000011100000000000",--7291
"001111001110000010000000000000000010",--7292
"111110010000001010010100000000000000",--7293
"111110001110000010000011100000000000",--7294
"001101001100000001100000000000000110",--7295
"011010001111000000000000000000000010",--7296
"011111001101000000010000000000101000",--7297
"000101000000000000000001110100010010",--7298
"011100001101000000000000000000100110",--7299
"000101000000000000000001110100010010",--7300
"111110001110001001110101000000000000",--7301
"001101001100000010000000000000000100",--7302
"001111010000000010110000000000000000",--7303
"111110010100001010110101000000000000",--7304
"111110010000001010000101100000000000",--7305
"001111010000000011000000000000000001",--7306
"111110010110001011000101100000000000",--7307
"111110010100000010110101000000000000",--7308
"111110010010001010010101100000000000",--7309
"001111010000000011000000000000000010",--7310
"111110010110001011000101100000000000",--7311
"111110010100000010110101000000000000",--7312
"001101001100000010000000000000000011",--7313
"011100010001000000000000000000000011",--7314
"101110010101111000000011100000000000",--7315
"011111001111000000110000000000010000",--7316
"000101000000000000000001110010100100",--7317
"111110010000001010010101100000000000",--7318
"001101001100000010000000000000001001",--7319
"001111010000000011000000000000000000",--7320
"111110010110001011000101100000000000",--7321
"111110010100000010110101000000000000",--7322
"111110010010001001110100100000000000",--7323
"001111010000000010110000000000000001",--7324
"111110010010001010110100100000000000",--7325
"111110010100000010010100100000000000",--7326
"111110001110001010000011100000000000",--7327
"001111010000000010000000000000000010",--7328
"111110001110001010000011100000000000",--7329
"111110010010000001110011100000000000",--7330
"011111001111000000110000000000000001",--7331
"111110001110010000010011100000000000",--7332
"001101001100000001100000000000000110",--7333
"011010001111000000000000000000000010",--7334
"011111001101000000010000000000000010",--7335
"000101000000000000000001110100010010",--7336
"010000001101000000000000000001101000",--7337
"001101000110000001100000000000000001",--7338
"010011001101000000000000000001011010",--7339
"001101001100000001100000000101101101",--7340
"001101001100000001110000000000000101",--7341
"001111001110000001110000000000000000",--7342
"111110001000010001110011100000000000",--7343
"001111001110000010000000000000000001",--7344
"111110001010010010000100000000000000",--7345
"001111001110000010010000000000000010",--7346
"111110001100010010010100100000000000",--7347
"001101001100000001110000000000000001",--7348
"011111001111000000010000000000010000",--7349
"101110001111111000000011100000000001",--7350
"001101001100000001110000000000000100",--7351
"001111001110000010100000000000000000",--7352
"010110010101000001110000000000001001",--7353
"101110010001111000000011100000000001",--7354
"001111001110000010000000000000000001",--7355
"010110010001000001110000000000000110",--7356
"101110010011111000000011100000000001",--7357
"001111001110000010000000000000000010",--7358
"010110010001000001110000000000000011",--7359
"001101001100000001100000000000000110",--7360
"011100001101000000000000000001010000",--7361
"000101000000000000000001110011111011",--7362
"001101001100000001100000000000000110",--7363
"011100001101000000000000000000110110",--7364
"000101000000000000000001110100010010",--7365
"011111001111000000100000000000001111",--7366
"001101001100000001110000000000000100",--7367
"001111001110000010100000000000000000",--7368
"111110010100001001110011100000000000",--7369
"001111001110000010100000000000000001",--7370
"111110010100001010000100000000000000",--7371
"111110001110000010000011100000000000",--7372
"001111001110000010000000000000000010",--7373
"111110010000001010010100000000000000",--7374
"111110001110000010000011100000000000",--7375
"001101001100000001100000000000000110",--7376
"011010001111000000000000000000000010",--7377
"011111001101000000010000000000101000",--7378
"000101000000000000000001110100010010",--7379
"011100001101000000000000000000100110",--7380
"000101000000000000000001110100010010",--7381
"111110001110001001110101000000000000",--7382
"001101001100000010000000000000000100",--7383
"001111010000000010110000000000000000",--7384
"111110010100001010110101000000000000",--7385
"111110010000001010000101100000000000",--7386
"001111010000000011000000000000000001",--7387
"111110010110001011000101100000000000",--7388
"111110010100000010110101000000000000",--7389
"111110010010001010010101100000000000",--7390
"001111010000000011000000000000000010",--7391
"111110010110001011000101100000000000",--7392
"111110010100000010110101000000000000",--7393
"001101001100000010000000000000000011",--7394
"011100010001000000000000000000000011",--7395
"101110010101111000000011100000000000",--7396
"011111001111000000110000000000010000",--7397
"000101000000000000000001110011110101",--7398
"111110010000001010010101100000000000",--7399
"001101001100000010000000000000001001",--7400
"001111010000000011000000000000000000",--7401
"111110010110001011000101100000000000",--7402
"111110010100000010110101000000000000",--7403
"111110010010001001110100100000000000",--7404
"001111010000000010110000000000000001",--7405
"111110010010001010110100100000000000",--7406
"111110010100000010010100100000000000",--7407
"111110001110001010000011100000000000",--7408
"001111010000000010000000000000000010",--7409
"111110001110001010000011100000000000",--7410
"111110010010000001110011100000000000",--7411
"011111001111000000110000000000000001",--7412
"111110001110010000010011100000000000",--7413
"001101001100000001100000000000000110",--7414
"011010001111000000000000000000000010",--7415
"011111001101000000010000000000000010",--7416
"000101000000000000000001110100010010",--7417
"010000001101000000000000000000010111",--7418
"101000000111111000000001000000000000",--7419
"101001000000000000010000000000000010",--7420
"101110001001111000000001100000000000",--7421
"101110001011111000000010000000000000",--7422
"101110001101111000000010100000000000",--7423
"001001111100000111111111111111110110",--7424
"101001111100010111100000000000001011",--7425
"000111000000000000000000011110001000",--7426
"101001111100000111100000000000001011",--7427
"001101111100000111111111111111110110",--7428
"010000000011000000000000000000001100",--7429
"001111111100000000111111111111110111",--7430
"001011000000000000110000000100101101",--7431
"001111111100000000111111111111111000",--7432
"001011000000000000110000000100101010",--7433
"001111111100000000111111111111111001",--7434
"001011000000000000110000000100101011",--7435
"001111111100000000111111111111111010",--7436
"001011000000000000110000000100101100",--7437
"001101111100000000011111111111111011",--7438
"001001000000000000010000000100101001",--7439
"001101111100000000011111111111111100",--7440
"001001000000000000010000000100101110",--7441
"001101111100000000011111111111111101",--7442
"101001000010000000010000000000000001",--7443
"001101111100000000101111111111111111",--7444
"001101111100000000110000000000000000",--7445
"000101000000000000000001011101010010",--7446
"001100000100000000010010000000000000",--7447
"010011001000000000001111100000000000",--7448
"001101001000000001000000000100110001",--7449
"001101001000000001010000000000000000",--7450
"001001111100000000110000000000000000",--7451
"001001111100000000101111111111111111",--7452
"001001111100000000011111111111111110",--7453
"010011001011000000000000000111010110",--7454
"001101001010000001100000000101101101",--7455
"001111000000000000110000000100010101",--7456
"001101001100000001110000000000000101",--7457
"001111001110000001000000000000000000",--7458
"111110000110010001000001100000000000",--7459
"001111000000000001000000000100010110",--7460
"001111001110000001010000000000000001",--7461
"111110001000010001010010000000000000",--7462
"001111000000000001010000000100010111",--7463
"001111001110000001100000000000000010",--7464
"111110001010010001100010100000000000",--7465
"001101001100000001110000000000000001",--7466
"011111001111000000010000000001010100",--7467
"001111000110000001100000000000000000",--7468
"010010001101000000000000000000011010",--7469
"001101001100000001110000000000000100",--7470
"001101001100000010000000000000000110",--7471
"011010001101000000000000000000000010",--7472
"101001000000000010010000000000000001",--7473
"000101000000000000000001110100110100",--7474
"101000000001111000000100100000000000",--7475
"001111001110000001100000000000000000",--7476
"011100010001000010010000000000000001",--7477
"101110001101111000000011000000000010",--7478
"111110001100010000110011000000000000",--7479
"001111000110000001110000000000000000",--7480
"111110001110011000000011100000000000",--7481
"111110001100001001110011000000000000",--7482
"001111000110000001110000000000000001",--7483
"111110001100001001110011100000000000",--7484
"111110001110000001000011100000000001",--7485
"001111001110000010000000000000000001",--7486
"010110010001000001110000000000001000",--7487
"001111000110000001110000000000000010",--7488
"111110001100001001110011100000000000",--7489
"111110001110000001010011100000000001",--7490
"001111001110000010000000000000000010",--7491
"010110010001000001110000000000000011",--7492
"001011000000000001100000000100101111",--7493
"101001000000000001100000000000000001",--7494
"000101000000000000000001111000011010",--7495
"001111000110000001100000000000000001",--7496
"010010001101000000000000000000011010",--7497
"001101001100000001110000000000000100",--7498
"001101001100000010000000000000000110",--7499
"011010001101000000000000000000000010",--7500
"101001000000000010010000000000000001",--7501
"000101000000000000000001110101010000",--7502
"101000000001111000000100100000000000",--7503
"001111001110000001100000000000000001",--7504
"011100010001000010010000000000000001",--7505
"101110001101111000000011000000000010",--7506
"111110001100010001000011000000000000",--7507
"001111000110000001110000000000000001",--7508
"111110001110011000000011100000000000",--7509
"111110001100001001110011000000000000",--7510
"001111000110000001110000000000000010",--7511
"111110001100001001110011100000000000",--7512
"111110001110000001010011100000000001",--7513
"001111001110000010000000000000000010",--7514
"010110010001000001110000000000001000",--7515
"001111000110000001110000000000000000",--7516
"111110001100001001110011100000000000",--7517
"111110001110000000110011100000000001",--7518
"001111001110000010000000000000000000",--7519
"010110010001000001110000000000000011",--7520
"001011000000000001100000000100101111",--7521
"101001000000000001100000000000000010",--7522
"000101000000000000000001111000011010",--7523
"001111000110000001100000000000000010",--7524
"010010001101000000000000000010101001",--7525
"001101001100000001110000000000000100",--7526
"001101001100000001100000000000000110",--7527
"011010001101000000000000000000000010",--7528
"101001000000000010000000000000000001",--7529
"000101000000000000000001110101101100",--7530
"101000000001111000000100000000000000",--7531
"001111001110000001100000000000000010",--7532
"011100001101000010000000000000000001",--7533
"101110001101111000000011000000000010",--7534
"111110001100010001010010100000000000",--7535
"001111000110000001100000000000000010",--7536
"111110001100011000000011000000000000",--7537
"111110001010001001100010100000000000",--7538
"001111000110000001100000000000000000",--7539
"111110001010001001100011000000000000",--7540
"111110001100000000110001100000000001",--7541
"001111001110000001100000000000000000",--7542
"010110001101000000110000000010010111",--7543
"001111000110000000110000000000000001",--7544
"111110001010001000110001100000000000",--7545
"111110000110000001000001100000000001",--7546
"001111001110000001000000000000000001",--7547
"010110001001000000110000000010010010",--7548
"001011000000000001010000000100101111",--7549
"101001000000000001100000000000000011",--7550
"000101000000000000000001111000011010",--7551
"011111001111000000100000000000011010",--7552
"001101001100000001100000000000000100",--7553
"001111000110000001100000000000000000",--7554
"001111001100000001110000000000000000",--7555
"111110001100001001110011000000000000",--7556
"001111000110000001110000000000000001",--7557
"001111001100000010000000000000000001",--7558
"111110001110001010000011100000000000",--7559
"111110001100000001110011000000000000",--7560
"001111000110000001110000000000000010",--7561
"001111001100000010000000000000000010",--7562
"111110001110001010000011100000000000",--7563
"111110001100000001110011000000000000",--7564
"010110001101000000000000000010000001",--7565
"001111001100000001110000000000000000",--7566
"111110001110001000110001100000000000",--7567
"001111001100000001110000000000000001",--7568
"111110001110001001000010000000000000",--7569
"111110000110000001000001100000000000",--7570
"001111001100000001000000000000000010",--7571
"111110001000001001010010000000000000",--7572
"111110000110000001000001100000000010",--7573
"111110001100011000000010000000000000",--7574
"111110000110001001000001100000000000",--7575
"001011000000000000110000000100101111",--7576
"101001000000000001100000000000000001",--7577
"000101000000000000000001111000011010",--7578
"001111000110000001100000000000000000",--7579
"001111000110000001110000000000000001",--7580
"001111000110000010000000000000000010",--7581
"111110001100001001100100100000000000",--7582
"001101001100000010000000000000000100",--7583
"001111010000000010100000000000000000",--7584
"111110010010001010100100100000000000",--7585
"111110001110001001110101000000000000",--7586
"001111010000000010110000000000000001",--7587
"111110010100001010110101000000000000",--7588
"111110010010000010100100100000000000",--7589
"111110010000001010000101000000000000",--7590
"001111010000000010110000000000000010",--7591
"111110010100001010110101000000000000",--7592
"111110010010000010100100100000000000",--7593
"001101001100000010010000000000000011",--7594
"011100010011000000000000000000000011",--7595
"101110010011111000000011000000000000",--7596
"011110010011000000000000000000001111",--7597
"000101000000000000000001111000001111",--7598
"111110001110001010000101000000000000",--7599
"001101001100000010100000000000001001",--7600
"001111010100000010110000000000000000",--7601
"111110010100001010110101000000000000",--7602
"111110010010000010100100100000000000",--7603
"111110010000001001100100000000000000",--7604
"001111010100000010100000000000000001",--7605
"111110010000001010100100000000000000",--7606
"111110010010000010000100000000000000",--7607
"111110001100001001110011000000000000",--7608
"001111010100000001110000000000000010",--7609
"111110001100001001110011000000000000",--7610
"111110010000000001100011000000000000",--7611
"010010001101000000000000000001010010",--7612
"001111000110000001110000000000000000",--7613
"001111000110000010000000000000000001",--7614
"001111000110000010010000000000000010",--7615
"111110001110001000110101000000000000",--7616
"001111010000000010110000000000000000",--7617
"111110010100001010110101000000000000",--7618
"111110010000001001000101100000000000",--7619
"001111010000000011000000000000000001",--7620
"111110010110001011000101100000000000",--7621
"111110010100000010110101000000000000",--7622
"111110010010001001010101100000000000",--7623
"001111010000000011000000000000000010",--7624
"111110010110001011000101100000000000",--7625
"111110010100000010110101000000000000",--7626
"011100010011000000000000000000000010",--7627
"101110010101111000000011100000000000",--7628
"000101000000000000000001110111100011",--7629
"111110010010001001000101100000000000",--7630
"111110010000001001010110000000000000",--7631
"111110010110000011000101100000000000",--7632
"001101001100000010100000000000001001",--7633
"001111010100000011000000000000000000",--7634
"111110010110001011000101100000000000",--7635
"111110001110001001010110000000000000",--7636
"111110010010001000110100100000000000",--7637
"111110011000000010010100100000000000",--7638
"001111010100000011000000000000000001",--7639
"111110010010001011000100100000000000",--7640
"111110010110000010010100100000000000",--7641
"111110001110001001000011100000000000",--7642
"111110010000001000110100000000000000",--7643
"111110001110000010000011100000000000",--7644
"001111010100000010000000000000000010",--7645
"111110001110001010000011100000000000",--7646
"111110010010000001110011100000000000",--7647
"101111000001110010000011111100000000",--7648
"111110001110001010000011100000000000",--7649
"111110010100000001110011100000000000",--7650
"111110000110001000110100000000000000",--7651
"001111010000000010010000000000000000",--7652
"111110010000001010010100000000000000",--7653
"111110001000001001000100100000000000",--7654
"001111010000000010100000000000000001",--7655
"111110010010001010100100100000000000",--7656
"111110010000000010010100000000000000",--7657
"111110001010001001010100100000000000",--7658
"001111010000000010100000000000000010",--7659
"111110010010001010100100100000000000",--7660
"111110010000000010010100000000000000",--7661
"011100010011000000000000000000000011",--7662
"101110010001111000000001100000000000",--7663
"011111001111000000110000000000010000",--7664
"000101000000000000000001111000000000",--7665
"111110001000001001010100100000000000",--7666
"001101001100000010000000000000001001",--7667
"001111010000000010100000000000000000",--7668
"111110010010001010100100100000000000",--7669
"111110010000000010010100000000000000",--7670
"111110001010001000110010100000000000",--7671
"001111010000000010010000000000000001",--7672
"111110001010001010010010100000000000",--7673
"111110010000000001010010100000000000",--7674
"111110000110001001000001100000000000",--7675
"001111010000000001000000000000000010",--7676
"111110000110001001000001100000000000",--7677
"111110001010000000110001100000000000",--7678
"011111001111000000110000000000000001",--7679
"111110000110010000010001100000000000",--7680
"111110001110001001110010000000000000",--7681
"111110001100001000110001100000000000",--7682
"111110001000010000110001100000000000",--7683
"010110000111000000000000000000001010",--7684
"111110000110100000000001100000000000",--7685
"001101001100000001100000000000000110",--7686
"011100001101000000000000000000000001",--7687
"101110000111111000000001100000000010",--7688
"111110000110010001110001100000000000",--7689
"111110001100011000000010000000000000",--7690
"111110000110001001000001100000000000",--7691
"001011000000000000110000000100101111",--7692
"101001000000000001100000000000000001",--7693
"000101000000000000000001111000011010",--7694
"001101001010000001010000000101101101",--7695
"001101001010000001010000000000000110",--7696
"010000001011000000000000000011100011",--7697
"101000001001111000000001000000000000",--7698
"101001000000000000010000000000000001",--7699
"001001111100000111111111111111111101",--7700
"101001111100010111100000000000000100",--7701
"000111000000000000000001011101010010",--7702
"101001111100000111100000000000000100",--7703
"001101111100000111111111111111111101",--7704
"000101000000000000000001111011110101",--7705
"001111000000000000110000000100101111",--7706
"001001111100000001001111111111111101",--7707
"010110000111000000000000000011010000",--7708
"001111000000000001000000000100101101",--7709
"010110001001000000110000000011001110",--7710
"101111001001110001000011110000100011",--7711
"101111001001100001001101011100001010",--7712
"111110000110000001000001100000000000",--7713
"001111000110000001000000000000000000",--7714
"111110001000001000110010000000000000",--7715
"001111000000000001010000000100010101",--7716
"111110001000000001010010000000000000",--7717
"001111000110000001010000000000000001",--7718
"111110001010001000110010100000000000",--7719
"001111000000000001100000000100010110",--7720
"111110001010000001100010100000000000",--7721
"001111000110000001100000000000000010",--7722
"111110001100001000110011000000000000",--7723
"001111000000000001110000000100010111",--7724
"111110001100000001110011000000000000",--7725
"001101001000000001110000000000000000",--7726
"001001111100000001101111111111111100",--7727
"001001111100000001011111111111111011",--7728
"001011111100000001101111111111111010",--7729
"001011111100000001011111111111111001",--7730
"001011111100000001001111111111111000",--7731
"001011111100000000111111111111110111",--7732
"010011001111000000000000000010101011",--7733
"001101001110000001110000000101101101",--7734
"001101001110000010000000000000000101",--7735
"001111010000000001110000000000000000",--7736
"111110001000010001110011100000000000",--7737
"001111010000000010000000000000000001",--7738
"111110001010010010000100000000000000",--7739
"001111010000000010010000000000000010",--7740
"111110001100010010010100100000000000",--7741
"001101001110000010000000000000000001",--7742
"011111010001000000010000000000010000",--7743
"101110001111111000000011100000000001",--7744
"001101001110000010000000000000000100",--7745
"001111010000000010100000000000000000",--7746
"010110010101000001110000000000001001",--7747
"101110010001111000000011100000000001",--7748
"001111010000000010000000000000000001",--7749
"010110010001000001110000000000000110",--7750
"101110010011111000000011100000000001",--7751
"001111010000000010000000000000000010",--7752
"010110010001000001110000000000000011",--7753
"001101001110000001110000000000000110",--7754
"011100001111000000000000000010100001",--7755
"000101000000000000000001111010000101",--7756
"001101001110000001110000000000000110",--7757
"011100001111000000000000000000110110",--7758
"000101000000000000000001111011101101",--7759
"011111010001000000100000000000001111",--7760
"001101001110000010000000000000000100",--7761
"001111010000000010100000000000000000",--7762
"111110010100001001110011100000000000",--7763
"001111010000000010100000000000000001",--7764
"111110010100001010000100000000000000",--7765
"111110001110000010000011100000000000",--7766
"001111010000000010000000000000000010",--7767
"111110010000001010010100000000000000",--7768
"111110001110000010000011100000000000",--7769
"001101001110000001110000000000000110",--7770
"011010001111000000000000000000000010",--7771
"011111001111000000010000000000101000",--7772
"000101000000000000000001111011101101",--7773
"011100001111000000000000000000100110",--7774
"000101000000000000000001111011101101",--7775
"111110001110001001110101000000000000",--7776
"001101001110000010010000000000000100",--7777
"001111010010000010110000000000000000",--7778
"111110010100001010110101000000000000",--7779
"111110010000001010000101100000000000",--7780
"001111010010000011000000000000000001",--7781
"111110010110001011000101100000000000",--7782
"111110010100000010110101000000000000",--7783
"111110010010001010010101100000000000",--7784
"001111010010000011000000000000000010",--7785
"111110010110001011000101100000000000",--7786
"111110010100000010110101000000000000",--7787
"001101001110000010010000000000000011",--7788
"011100010011000000000000000000000011",--7789
"101110010101111000000011100000000000",--7790
"011111010001000000110000000000010000",--7791
"000101000000000000000001111001111111",--7792
"111110010000001010010101100000000000",--7793
"001101001110000010010000000000001001",--7794
"001111010010000011000000000000000000",--7795
"111110010110001011000101100000000000",--7796
"111110010100000010110101000000000000",--7797
"111110010010001001110100100000000000",--7798
"001111010010000010110000000000000001",--7799
"111110010010001010110100100000000000",--7800
"111110010100000010010100100000000000",--7801
"111110001110001010000011100000000000",--7802
"001111010010000010000000000000000010",--7803
"111110001110001010000011100000000000",--7804
"111110010010000001110011100000000000",--7805
"011111010001000000110000000000000001",--7806
"111110001110010000010011100000000000",--7807
"001101001110000001110000000000000110",--7808
"011010001111000000000000000000000010",--7809
"011111001111000000010000000000000010",--7810
"000101000000000000000001111011101101",--7811
"010000001111000000000000000001101000",--7812
"001101001000000001110000000000000001",--7813
"010011001111000000000000000001011010",--7814
"001101001110000001110000000101101101",--7815
"001101001110000010000000000000000101",--7816
"001111010000000001110000000000000000",--7817
"111110001000010001110011100000000000",--7818
"001111010000000010000000000000000001",--7819
"111110001010010010000100000000000000",--7820
"001111010000000010010000000000000010",--7821
"111110001100010010010100100000000000",--7822
"001101001110000010000000000000000001",--7823
"011111010001000000010000000000010000",--7824
"101110001111111000000011100000000001",--7825
"001101001110000010000000000000000100",--7826
"001111010000000010100000000000000000",--7827
"010110010101000001110000000000001001",--7828
"101110010001111000000011100000000001",--7829
"001111010000000010000000000000000001",--7830
"010110010001000001110000000000000110",--7831
"101110010011111000000011100000000001",--7832
"001111010000000010000000000000000010",--7833
"010110010001000001110000000000000011",--7834
"001101001110000001110000000000000110",--7835
"011100001111000000000000000001010000",--7836
"000101000000000000000001111011010110",--7837
"001101001110000001110000000000000110",--7838
"011100001111000000000000000000110110",--7839
"000101000000000000000001111011101101",--7840
"011111010001000000100000000000001111",--7841
"001101001110000010000000000000000100",--7842
"001111010000000010100000000000000000",--7843
"111110010100001001110011100000000000",--7844
"001111010000000010100000000000000001",--7845
"111110010100001010000100000000000000",--7846
"111110001110000010000011100000000000",--7847
"001111010000000010000000000000000010",--7848
"111110010000001010010100000000000000",--7849
"111110001110000010000011100000000000",--7850
"001101001110000001110000000000000110",--7851
"011010001111000000000000000000000010",--7852
"011111001111000000010000000000101000",--7853
"000101000000000000000001111011101101",--7854
"011100001111000000000000000000100110",--7855
"000101000000000000000001111011101101",--7856
"111110001110001001110101000000000000",--7857
"001101001110000010010000000000000100",--7858
"001111010010000010110000000000000000",--7859
"111110010100001010110101000000000000",--7860
"111110010000001010000101100000000000",--7861
"001111010010000011000000000000000001",--7862
"111110010110001011000101100000000000",--7863
"111110010100000010110101000000000000",--7864
"111110010010001010010101100000000000",--7865
"001111010010000011000000000000000010",--7866
"111110010110001011000101100000000000",--7867
"111110010100000010110101000000000000",--7868
"001101001110000010010000000000000011",--7869
"011100010011000000000000000000000011",--7870
"101110010101111000000011100000000000",--7871
"011111010001000000110000000000010000",--7872
"000101000000000000000001111011010000",--7873
"111110010000001010010101100000000000",--7874
"001101001110000010010000000000001001",--7875
"001111010010000011000000000000000000",--7876
"111110010110001011000101100000000000",--7877
"111110010100000010110101000000000000",--7878
"111110010010001001110100100000000000",--7879
"001111010010000010110000000000000001",--7880
"111110010010001010110100100000000000",--7881
"111110010100000010010100100000000000",--7882
"111110001110001010000011100000000000",--7883
"001111010010000010000000000000000010",--7884
"111110001110001010000011100000000000",--7885
"111110010010000001110011100000000000",--7886
"011111010001000000110000000000000001",--7887
"111110001110010000010011100000000000",--7888
"001101001110000001110000000000000110",--7889
"011010001111000000000000000000000010",--7890
"011111001111000000010000000000000010",--7891
"000101000000000000000001111011101101",--7892
"010000001111000000000000000000010111",--7893
"101000001001111000000001000000000000",--7894
"101001000000000000010000000000000010",--7895
"101110001001111000000001100000000000",--7896
"101110001011111000000010000000000000",--7897
"101110001101111000000010100000000000",--7898
"001001111100000111111111111111110110",--7899
"101001111100010111100000000000001011",--7900
"000111000000000000000000011110001000",--7901
"101001111100000111100000000000001011",--7902
"001101111100000111111111111111110110",--7903
"010000000011000000000000000000001100",--7904
"001111111100000000111111111111110111",--7905
"001011000000000000110000000100101101",--7906
"001111111100000000111111111111111000",--7907
"001011000000000000110000000100101010",--7908
"001111111100000000111111111111111001",--7909
"001011000000000000110000000100101011",--7910
"001111111100000000111111111111111010",--7911
"001011000000000000110000000100101100",--7912
"001101111100000000011111111111111011",--7913
"001001000000000000010000000100101001",--7914
"001101111100000000011111111111111100",--7915
"001001000000000000010000000100101110",--7916
"101001000000000000010000000000000001",--7917
"001101111100000000101111111111111101",--7918
"001101111100000000110000000000000000",--7919
"001001111100000111111111111111111100",--7920
"101001111100010111100000000000000101",--7921
"000111000000000000000001011101010010",--7922
"101001111100000111100000000000000101",--7923
"001101111100000111111111111111111100",--7924
"001101111100000000011111111111111110",--7925
"101001000010000000010000000000000001",--7926
"001101111100000000111111111111111111",--7927
"001100000110000000010001000000000000",--7928
"010011000100000000001111100000000000",--7929
"001101000100000000100000000100110001",--7930
"001101111100000000110000000000000000",--7931
"001001111100000000011111111111111101",--7932
"101000000001111000000000100000000000",--7933
"001001111100000111111111111111111100",--7934
"101001111100010111100000000000000101",--7935
"000111000000000000000001011101010010",--7936
"101001111100000111100000000000000101",--7937
"001101111100000111111111111111111100",--7938
"001101111100000000011111111111111101",--7939
"101001000010000000010000000000000001",--7940
"001101111100000000111111111111111111",--7941
"001100000110000000010001000000000000",--7942
"010011000100000000001111100000000000",--7943
"001101000100000000100000000100110001",--7944
"001101000100000001000000000000000000",--7945
"001001111100000000011111111111111100",--7946
"010011001001000000000000000100110111",--7947
"001101001000000001010000000101101101",--7948
"001111000000000000110000000100010101",--7949
"001101001010000001100000000000000101",--7950
"001111001100000001000000000000000000",--7951
"111110000110010001000001100000000000",--7952
"001111000000000001000000000100010110",--7953
"001111001100000001010000000000000001",--7954
"111110001000010001010010000000000000",--7955
"001111000000000001010000000100010111",--7956
"001111001100000001100000000000000010",--7957
"111110001010010001100010100000000000",--7958
"001101001010000001100000000000000001",--7959
"011111001101000000010000000001010101",--7960
"001101111100000001100000000000000000",--7961
"001111001100000001100000000000000000",--7962
"010010001101000000000000000000011010",--7963
"001101001010000001110000000000000100",--7964
"001101001010000010000000000000000110",--7965
"011010001101000000000000000000000010",--7966
"101001000000000010010000000000000001",--7967
"000101000000000000000001111100100010",--7968
"101000000001111000000100100000000000",--7969
"001111001110000001100000000000000000",--7970
"011100010001000010010000000000000001",--7971
"101110001101111000000011000000000010",--7972
"111110001100010000110011000000000000",--7973
"001111001100000001110000000000000000",--7974
"111110001110011000000011100000000000",--7975
"111110001100001001110011000000000000",--7976
"001111001100000001110000000000000001",--7977
"111110001100001001110011100000000000",--7978
"111110001110000001000011100000000001",--7979
"001111001110000010000000000000000001",--7980
"010110010001000001110000000000001000",--7981
"001111001100000001110000000000000010",--7982
"111110001100001001110011100000000000",--7983
"111110001110000001010011100000000001",--7984
"001111001110000010000000000000000010",--7985
"010110010001000001110000000000000011",--7986
"001011000000000001100000000100101111",--7987
"101001000000000001010000000000000001",--7988
"000101000000000000000010000000001010",--7989
"001111001100000001100000000000000001",--7990
"010010001101000000000000000000011010",--7991
"001101001010000001110000000000000100",--7992
"001101001010000010000000000000000110",--7993
"011010001101000000000000000000000010",--7994
"101001000000000010010000000000000001",--7995
"000101000000000000000001111100111110",--7996
"101000000001111000000100100000000000",--7997
"001111001110000001100000000000000001",--7998
"011100010001000010010000000000000001",--7999
"101110001101111000000011000000000010",--8000
"111110001100010001000011000000000000",--8001
"001111001100000001110000000000000001",--8002
"111110001110011000000011100000000000",--8003
"111110001100001001110011000000000000",--8004
"001111001100000001110000000000000010",--8005
"111110001100001001110011100000000000",--8006
"111110001110000001010011100000000001",--8007
"001111001110000010000000000000000010",--8008
"010110010001000001110000000000001000",--8009
"001111001100000001110000000000000000",--8010
"111110001100001001110011100000000000",--8011
"111110001110000000110011100000000001",--8012
"001111001110000010000000000000000000",--8013
"010110010001000001110000000000000011",--8014
"001011000000000001100000000100101111",--8015
"101001000000000001010000000000000010",--8016
"000101000000000000000010000000001010",--8017
"001111001100000001100000000000000010",--8018
"010010001101000000000000000010101011",--8019
"001101001010000001110000000000000100",--8020
"001101001010000001010000000000000110",--8021
"011010001101000000000000000000000010",--8022
"101001000000000010000000000000000001",--8023
"000101000000000000000001111101011010",--8024
"101000000001111000000100000000000000",--8025
"001111001110000001100000000000000010",--8026
"011100001011000010000000000000000001",--8027
"101110001101111000000011000000000010",--8028
"111110001100010001010010100000000000",--8029
"001111001100000001100000000000000010",--8030
"111110001100011000000011000000000000",--8031
"111110001010001001100010100000000000",--8032
"001111001100000001100000000000000000",--8033
"111110001010001001100011000000000000",--8034
"111110001100000000110001100000000001",--8035
"001111001110000001100000000000000000",--8036
"010110001101000000110000000010011001",--8037
"001111001100000000110000000000000001",--8038
"111110001010001000110001100000000000",--8039
"111110000110000001000001100000000001",--8040
"001111001110000001000000000000000001",--8041
"010110001001000000110000000010010100",--8042
"001011000000000001010000000100101111",--8043
"101001000000000001010000000000000011",--8044
"000101000000000000000010000000001010",--8045
"011111001101000000100000000000011011",--8046
"001101001010000001010000000000000100",--8047
"001101111100000001100000000000000000",--8048
"001111001100000001100000000000000000",--8049
"001111001010000001110000000000000000",--8050
"111110001100001001110011000000000000",--8051
"001111001100000001110000000000000001",--8052
"001111001010000010000000000000000001",--8053
"111110001110001010000011100000000000",--8054
"111110001100000001110011000000000000",--8055
"001111001100000001110000000000000010",--8056
"001111001010000010000000000000000010",--8057
"111110001110001010000011100000000000",--8058
"111110001100000001110011000000000000",--8059
"010110001101000000000000000010000010",--8060
"001111001010000001110000000000000000",--8061
"111110001110001000110001100000000000",--8062
"001111001010000001110000000000000001",--8063
"111110001110001001000010000000000000",--8064
"111110000110000001000001100000000000",--8065
"001111001010000001000000000000000010",--8066
"111110001000001001010010000000000000",--8067
"111110000110000001000001100000000010",--8068
"111110001100011000000010000000000000",--8069
"111110000110001001000001100000000000",--8070
"001011000000000000110000000100101111",--8071
"101001000000000001010000000000000001",--8072
"000101000000000000000010000000001010",--8073
"001101111100000001110000000000000000",--8074
"001111001110000001100000000000000000",--8075
"001111001110000001110000000000000001",--8076
"001111001110000010000000000000000010",--8077
"111110001100001001100100100000000000",--8078
"001101001010000010000000000000000100",--8079
"001111010000000010100000000000000000",--8080
"111110010010001010100100100000000000",--8081
"111110001110001001110101000000000000",--8082
"001111010000000010110000000000000001",--8083
"111110010100001010110101000000000000",--8084
"111110010010000010100100100000000000",--8085
"111110010000001010000101000000000000",--8086
"001111010000000010110000000000000010",--8087
"111110010100001010110101000000000000",--8088
"111110010010000010100100100000000000",--8089
"001101001010000010010000000000000011",--8090
"011100010011000000000000000000000011",--8091
"101110010011111000000011000000000000",--8092
"011110010011000000000000000000001111",--8093
"000101000000000000000001111111111111",--8094
"111110001110001010000101000000000000",--8095
"001101001010000010100000000000001001",--8096
"001111010100000010110000000000000000",--8097
"111110010100001010110101000000000000",--8098
"111110010010000010100100100000000000",--8099
"111110010000001001100100000000000000",--8100
"001111010100000010100000000000000001",--8101
"111110010000001010100100000000000000",--8102
"111110010010000010000100000000000000",--8103
"111110001100001001110011000000000000",--8104
"001111010100000001110000000000000010",--8105
"111110001100001001110011000000000000",--8106
"111110010000000001100011000000000000",--8107
"010010001101000000000000000001010010",--8108
"001111001110000001110000000000000000",--8109
"001111001110000010000000000000000001",--8110
"001111001110000010010000000000000010",--8111
"111110001110001000110101000000000000",--8112
"001111010000000010110000000000000000",--8113
"111110010100001010110101000000000000",--8114
"111110010000001001000101100000000000",--8115
"001111010000000011000000000000000001",--8116
"111110010110001011000101100000000000",--8117
"111110010100000010110101000000000000",--8118
"111110010010001001010101100000000000",--8119
"001111010000000011000000000000000010",--8120
"111110010110001011000101100000000000",--8121
"111110010100000010110101000000000000",--8122
"011100010011000000000000000000000010",--8123
"101110010101111000000011100000000000",--8124
"000101000000000000000001111111010011",--8125
"111110010010001001000101100000000000",--8126
"111110010000001001010110000000000000",--8127
"111110010110000011000101100000000000",--8128
"001101001010000010100000000000001001",--8129
"001111010100000011000000000000000000",--8130
"111110010110001011000101100000000000",--8131
"111110001110001001010110000000000000",--8132
"111110010010001000110100100000000000",--8133
"111110011000000010010100100000000000",--8134
"001111010100000011000000000000000001",--8135
"111110010010001011000100100000000000",--8136
"111110010110000010010100100000000000",--8137
"111110001110001001000011100000000000",--8138
"111110010000001000110100000000000000",--8139
"111110001110000010000011100000000000",--8140
"001111010100000010000000000000000010",--8141
"111110001110001010000011100000000000",--8142
"111110010010000001110011100000000000",--8143
"101111000001110010000011111100000000",--8144
"111110001110001010000011100000000000",--8145
"111110010100000001110011100000000000",--8146
"111110000110001000110100000000000000",--8147
"001111010000000010010000000000000000",--8148
"111110010000001010010100000000000000",--8149
"111110001000001001000100100000000000",--8150
"001111010000000010100000000000000001",--8151
"111110010010001010100100100000000000",--8152
"111110010000000010010100000000000000",--8153
"111110001010001001010100100000000000",--8154
"001111010000000010100000000000000010",--8155
"111110010010001010100100100000000000",--8156
"111110010000000010010100000000000000",--8157
"011100010011000000000000000000000011",--8158
"101110010001111000000001100000000000",--8159
"011111001101000000110000000000010000",--8160
"000101000000000000000001111111110000",--8161
"111110001000001001010100100000000000",--8162
"001101001010000010000000000000001001",--8163
"001111010000000010100000000000000000",--8164
"111110010010001010100100100000000000",--8165
"111110010000000010010100000000000000",--8166
"111110001010001000110010100000000000",--8167
"001111010000000010010000000000000001",--8168
"111110001010001010010010100000000000",--8169
"111110010000000001010010100000000000",--8170
"111110000110001001000001100000000000",--8171
"001111010000000001000000000000000010",--8172
"111110000110001001000001100000000000",--8173
"111110001010000000110001100000000000",--8174
"011111001101000000110000000000000001",--8175
"111110000110010000010001100000000000",--8176
"111110001110001001110010000000000000",--8177
"111110001100001000110001100000000000",--8178
"111110001000010000110001100000000000",--8179
"010110000111000000000000000000001010",--8180
"111110000110100000000001100000000000",--8181
"001101001010000001010000000000000110",--8182
"011100001011000000000000000000000001",--8183
"101110000111111000000001100000000010",--8184
"111110000110010001110001100000000000",--8185
"111110001100011000000010000000000000",--8186
"111110000110001001000001100000000000",--8187
"001011000000000000110000000100101111",--8188
"101001000000000001010000000000000001",--8189
"000101000000000000000010000000001010",--8190
"001101001000000001000000000101101101",--8191
"001101001000000001000000000000000110",--8192
"010000001001000000000000000001000001",--8193
"001101111100000000110000000000000000",--8194
"101001000000000000010000000000000001",--8195
"001001111100000111111111111111111011",--8196
"101001111100010111100000000000000110",--8197
"000111000000000000000001011101010010",--8198
"101001111100000111100000000000000110",--8199
"001101111100000111111111111111111011",--8200
"000101000000000000000010000001000011",--8201
"001111000000000000110000000100101111",--8202
"001001111100000000101111111111111011",--8203
"010110000111000000000000000000101110",--8204
"001111000000000001000000000100101101",--8205
"010110001001000000110000000000101100",--8206
"101111001001110001000011110000100011",--8207
"101111001001100001001101011100001010",--8208
"111110000110000001000001100000000000",--8209
"001101111100000001100000000000000000",--8210
"001111001100000001000000000000000000",--8211
"111110001000001000110010000000000000",--8212
"001111000000000001010000000100010101",--8213
"111110001000000001010010000000000000",--8214
"001111001100000001010000000000000001",--8215
"111110001010001000110010100000000000",--8216
"001111000000000001100000000100010110",--8217
"111110001010000001100010100000000000",--8218
"001111001100000001100000000000000010",--8219
"111110001100001000110011000000000000",--8220
"001111000000000001110000000100010111",--8221
"111110001100000001110011000000000000",--8222
"001001111100000001011111111111111010",--8223
"001001111100000001001111111111111001",--8224
"001011111100000001101111111111111000",--8225
"001011111100000001011111111111110111",--8226
"001011111100000001001111111111110110",--8227
"001011111100000000111111111111110101",--8228
"101000000001111000000000100000000000",--8229
"101110001001111000000001100000000000",--8230
"101110001011111000000010000000000000",--8231
"101110001101111000000010100000000000",--8232
"001001111100000111111111111111110100",--8233
"101001111100010111100000000000001101",--8234
"000111000000000000000000011110001000",--8235
"101001111100000111100000000000001101",--8236
"001101111100000111111111111111110100",--8237
"010000000011000000000000000000001100",--8238
"001111111100000000111111111111110101",--8239
"001011000000000000110000000100101101",--8240
"001111111100000000111111111111110110",--8241
"001011000000000000110000000100101010",--8242
"001111111100000000111111111111110111",--8243
"001011000000000000110000000100101011",--8244
"001111111100000000111111111111111000",--8245
"001011000000000000110000000100101100",--8246
"001101111100000000011111111111111001",--8247
"001001000000000000010000000100101001",--8248
"001101111100000000011111111111111010",--8249
"001001000000000000010000000100101110",--8250
"101001000000000000010000000000000001",--8251
"001101111100000000101111111111111011",--8252
"001101111100000000110000000000000000",--8253
"001001111100000111111111111111111010",--8254
"101001111100010111100000000000000111",--8255
"000111000000000000000001011101010010",--8256
"101001111100000111100000000000000111",--8257
"001101111100000111111111111111111010",--8258
"001101111100000000011111111111111100",--8259
"101001000010000000010000000000000001",--8260
"001101111100000000111111111111111111",--8261
"001100000110000000010001000000000000",--8262
"010011000100000000001111100000000000",--8263
"001101000100000000100000000100110001",--8264
"001101111100000000110000000000000000",--8265
"001001111100000000011111111111111011",--8266
"101000000001111000000000100000000000",--8267
"001001111100000111111111111111111010",--8268
"101001111100010111100000000000000111",--8269
"000111000000000000000001011101010010",--8270
"101001111100000111100000000000000111",--8271
"001101111100000111111111111111111010",--8272
"001101111100000000011111111111111011",--8273
"101001000010000000010000000000000001",--8274
"001101111100000000101111111111111111",--8275
"001101111100000000110000000000000000",--8276
"000101000000000000000001110100010111",--8277
"001100000100000000010010000000000000",--8278
"001101001000000001010000000000000000",--8279
"010011001010000000001111100000000000",--8280
"001001111100000000110000000000000000",--8281
"001001111100000000101111111111111111",--8282
"001001111100000000011111111111111110",--8283
"011111001011011000110000000101011001",--8284
"001101001000000001010000000000000001",--8285
"010011001011000000000000001110011100",--8286
"001101001010000000100000000100110001",--8287
"001001111100000001001111111111111101",--8288
"101000000001111000000000100000000000",--8289
"001001111100000111111111111111111100",--8290
"101001111100010111100000000000000101",--8291
"000111000000000000000001011101010010",--8292
"101001111100000111100000000000000101",--8293
"001101111100000111111111111111111100",--8294
"001101111100000000011111111111111101",--8295
"001101000010000000100000000000000010",--8296
"010011000101000000000000001110010001",--8297
"001101000100000000100000000100110001",--8298
"001101000100000000110000000000000000",--8299
"010011000111000000000000000100110111",--8300
"001101000110000001000000000101101101",--8301
"001111000000000000110000000100010101",--8302
"001101001000000001010000000000000101",--8303
"001111001010000001000000000000000000",--8304
"111110000110010001000001100000000000",--8305
"001111000000000001000000000100010110",--8306
"001111001010000001010000000000000001",--8307
"111110001000010001010010000000000000",--8308
"001111000000000001010000000100010111",--8309
"001111001010000001100000000000000010",--8310
"111110001010010001100010100000000000",--8311
"001101001000000001010000000000000001",--8312
"011111001011000000010000000001010101",--8313
"001101111100000001010000000000000000",--8314
"001111001010000001100000000000000000",--8315
"010010001101000000000000000000011010",--8316
"001101001000000001100000000000000100",--8317
"001101001000000001110000000000000110",--8318
"011010001101000000000000000000000010",--8319
"101001000000000010000000000000000001",--8320
"000101000000000000000010000010000011",--8321
"101000000001111000000100000000000000",--8322
"001111001100000001100000000000000000",--8323
"011100001111000010000000000000000001",--8324
"101110001101111000000011000000000010",--8325
"111110001100010000110011000000000000",--8326
"001111001010000001110000000000000000",--8327
"111110001110011000000011100000000000",--8328
"111110001100001001110011000000000000",--8329
"001111001010000001110000000000000001",--8330
"111110001100001001110011100000000000",--8331
"111110001110000001000011100000000001",--8332
"001111001100000010000000000000000001",--8333
"010110010001000001110000000000001000",--8334
"001111001010000001110000000000000010",--8335
"111110001100001001110011100000000000",--8336
"111110001110000001010011100000000001",--8337
"001111001100000010000000000000000010",--8338
"010110010001000001110000000000000011",--8339
"001011000000000001100000000100101111",--8340
"101001000000000001000000000000000001",--8341
"000101000000000000000010000101101011",--8342
"001111001010000001100000000000000001",--8343
"010010001101000000000000000000011010",--8344
"001101001000000001100000000000000100",--8345
"001101001000000001110000000000000110",--8346
"011010001101000000000000000000000010",--8347
"101001000000000010000000000000000001",--8348
"000101000000000000000010000010011111",--8349
"101000000001111000000100000000000000",--8350
"001111001100000001100000000000000001",--8351
"011100001111000010000000000000000001",--8352
"101110001101111000000011000000000010",--8353
"111110001100010001000011000000000000",--8354
"001111001010000001110000000000000001",--8355
"111110001110011000000011100000000000",--8356
"111110001100001001110011000000000000",--8357
"001111001010000001110000000000000010",--8358
"111110001100001001110011100000000000",--8359
"111110001110000001010011100000000001",--8360
"001111001100000010000000000000000010",--8361
"010110010001000001110000000000001000",--8362
"001111001010000001110000000000000000",--8363
"111110001100001001110011100000000000",--8364
"111110001110000000110011100000000001",--8365
"001111001100000010000000000000000000",--8366
"010110010001000001110000000000000011",--8367
"001011000000000001100000000100101111",--8368
"101001000000000001000000000000000010",--8369
"000101000000000000000010000101101011",--8370
"001111001010000001100000000000000010",--8371
"010010001101000000000000000010101011",--8372
"001101001000000001100000000000000100",--8373
"001101001000000001000000000000000110",--8374
"011010001101000000000000000000000010",--8375
"101001000000000001110000000000000001",--8376
"000101000000000000000010000010111011",--8377
"101000000001111000000011100000000000",--8378
"001111001100000001100000000000000010",--8379
"011100001001000001110000000000000001",--8380
"101110001101111000000011000000000010",--8381
"111110001100010001010010100000000000",--8382
"001111001010000001100000000000000010",--8383
"111110001100011000000011000000000000",--8384
"111110001010001001100010100000000000",--8385
"001111001010000001100000000000000000",--8386
"111110001010001001100011000000000000",--8387
"111110001100000000110001100000000001",--8388
"001111001100000001100000000000000000",--8389
"010110001101000000110000000010011001",--8390
"001111001010000000110000000000000001",--8391
"111110001010001000110001100000000000",--8392
"111110000110000001000001100000000001",--8393
"001111001100000001000000000000000001",--8394
"010110001001000000110000000010010100",--8395
"001011000000000001010000000100101111",--8396
"101001000000000001000000000000000011",--8397
"000101000000000000000010000101101011",--8398
"011111001011000000100000000000011011",--8399
"001101001000000001000000000000000100",--8400
"001101111100000001010000000000000000",--8401
"001111001010000001100000000000000000",--8402
"001111001000000001110000000000000000",--8403
"111110001100001001110011000000000000",--8404
"001111001010000001110000000000000001",--8405
"001111001000000010000000000000000001",--8406
"111110001110001010000011100000000000",--8407
"111110001100000001110011000000000000",--8408
"001111001010000001110000000000000010",--8409
"001111001000000010000000000000000010",--8410
"111110001110001010000011100000000000",--8411
"111110001100000001110011000000000000",--8412
"010110001101000000000000000010000010",--8413
"001111001000000001110000000000000000",--8414
"111110001110001000110001100000000000",--8415
"001111001000000001110000000000000001",--8416
"111110001110001001000010000000000000",--8417
"111110000110000001000001100000000000",--8418
"001111001000000001000000000000000010",--8419
"111110001000001001010010000000000000",--8420
"111110000110000001000001100000000010",--8421
"111110001100011000000010000000000000",--8422
"111110000110001001000001100000000000",--8423
"001011000000000000110000000100101111",--8424
"101001000000000001000000000000000001",--8425
"000101000000000000000010000101101011",--8426
"001101111100000001100000000000000000",--8427
"001111001100000001100000000000000000",--8428
"001111001100000001110000000000000001",--8429
"001111001100000010000000000000000010",--8430
"111110001100001001100100100000000000",--8431
"001101001000000001110000000000000100",--8432
"001111001110000010100000000000000000",--8433
"111110010010001010100100100000000000",--8434
"111110001110001001110101000000000000",--8435
"001111001110000010110000000000000001",--8436
"111110010100001010110101000000000000",--8437
"111110010010000010100100100000000000",--8438
"111110010000001010000101000000000000",--8439
"001111001110000010110000000000000010",--8440
"111110010100001010110101000000000000",--8441
"111110010010000010100100100000000000",--8442
"001101001000000010000000000000000011",--8443
"011100010001000000000000000000000011",--8444
"101110010011111000000011000000000000",--8445
"011110010011000000000000000000001111",--8446
"000101000000000000000010000101100000",--8447
"111110001110001010000101000000000000",--8448
"001101001000000010010000000000001001",--8449
"001111010010000010110000000000000000",--8450
"111110010100001010110101000000000000",--8451
"111110010010000010100100100000000000",--8452
"111110010000001001100100000000000000",--8453
"001111010010000010100000000000000001",--8454
"111110010000001010100100000000000000",--8455
"111110010010000010000100000000000000",--8456
"111110001100001001110011000000000000",--8457
"001111010010000001110000000000000010",--8458
"111110001100001001110011000000000000",--8459
"111110010000000001100011000000000000",--8460
"010010001101000000000000000001010010",--8461
"001111001100000001110000000000000000",--8462
"001111001100000010000000000000000001",--8463
"001111001100000010010000000000000010",--8464
"111110001110001000110101000000000000",--8465
"001111001110000010110000000000000000",--8466
"111110010100001010110101000000000000",--8467
"111110010000001001000101100000000000",--8468
"001111001110000011000000000000000001",--8469
"111110010110001011000101100000000000",--8470
"111110010100000010110101000000000000",--8471
"111110010010001001010101100000000000",--8472
"001111001110000011000000000000000010",--8473
"111110010110001011000101100000000000",--8474
"111110010100000010110101000000000000",--8475
"011100010001000000000000000000000010",--8476
"101110010101111000000011100000000000",--8477
"000101000000000000000010000100110100",--8478
"111110010010001001000101100000000000",--8479
"111110010000001001010110000000000000",--8480
"111110010110000011000101100000000000",--8481
"001101001000000010010000000000001001",--8482
"001111010010000011000000000000000000",--8483
"111110010110001011000101100000000000",--8484
"111110001110001001010110000000000000",--8485
"111110010010001000110100100000000000",--8486
"111110011000000010010100100000000000",--8487
"001111010010000011000000000000000001",--8488
"111110010010001011000100100000000000",--8489
"111110010110000010010100100000000000",--8490
"111110001110001001000011100000000000",--8491
"111110010000001000110100000000000000",--8492
"111110001110000010000011100000000000",--8493
"001111010010000010000000000000000010",--8494
"111110001110001010000011100000000000",--8495
"111110010010000001110011100000000000",--8496
"101111000001110010000011111100000000",--8497
"111110001110001010000011100000000000",--8498
"111110010100000001110011100000000000",--8499
"111110000110001000110100000000000000",--8500
"001111001110000010010000000000000000",--8501
"111110010000001010010100000000000000",--8502
"111110001000001001000100100000000000",--8503
"001111001110000010100000000000000001",--8504
"111110010010001010100100100000000000",--8505
"111110010000000010010100000000000000",--8506
"111110001010001001010100100000000000",--8507
"001111001110000010100000000000000010",--8508
"111110010010001010100100100000000000",--8509
"111110010000000010010100000000000000",--8510
"011100010001000000000000000000000011",--8511
"101110010001111000000001100000000000",--8512
"011111001011000000110000000000010000",--8513
"000101000000000000000010000101010001",--8514
"111110001000001001010100100000000000",--8515
"001101001000000001110000000000001001",--8516
"001111001110000010100000000000000000",--8517
"111110010010001010100100100000000000",--8518
"111110010000000010010100000000000000",--8519
"111110001010001000110010100000000000",--8520
"001111001110000010010000000000000001",--8521
"111110001010001010010010100000000000",--8522
"111110010000000001010010100000000000",--8523
"111110000110001001000001100000000000",--8524
"001111001110000001000000000000000010",--8525
"111110000110001001000001100000000000",--8526
"111110001010000000110001100000000000",--8527
"011111001011000000110000000000000001",--8528
"111110000110010000010001100000000000",--8529
"111110001110001001110010000000000000",--8530
"111110001100001000110001100000000000",--8531
"111110001000010000110001100000000000",--8532
"010110000111000000000000000000001010",--8533
"111110000110100000000001100000000000",--8534
"001101001000000001000000000000000110",--8535
"011100001001000000000000000000000001",--8536
"101110000111111000000001100000000010",--8537
"111110000110010001110001100000000000",--8538
"111110001100011000000010000000000000",--8539
"111110000110001001000001100000000000",--8540
"001011000000000000110000000100101111",--8541
"101001000000000001000000000000000001",--8542
"000101000000000000000010000101101011",--8543
"001101000110000000110000000101101101",--8544
"001101000110000000110000000000000110",--8545
"010000000111000000000000000001000001",--8546
"001101111100000000110000000000000000",--8547
"101001000000000000010000000000000001",--8548
"001001111100000111111111111111111100",--8549
"101001111100010111100000000000000101",--8550
"000111000000000000000001011101010010",--8551
"101001111100000111100000000000000101",--8552
"001101111100000111111111111111111100",--8553
"000101000000000000000010000110100100",--8554
"001111000000000000110000000100101111",--8555
"001001111100000000101111111111111100",--8556
"010110000111000000000000000000101110",--8557
"001111000000000001000000000100101101",--8558
"010110001001000000110000000000101100",--8559
"101111001001110001000011110000100011",--8560
"101111001001100001001101011100001010",--8561
"111110000110000001000001100000000000",--8562
"001101111100000001010000000000000000",--8563
"001111001010000001000000000000000000",--8564
"111110001000001000110010000000000000",--8565
"001111000000000001010000000100010101",--8566
"111110001000000001010010000000000000",--8567
"001111001010000001010000000000000001",--8568
"111110001010001000110010100000000000",--8569
"001111000000000001100000000100010110",--8570
"111110001010000001100010100000000000",--8571
"001111001010000001100000000000000010",--8572
"111110001100001000110011000000000000",--8573
"001111000000000001110000000100010111",--8574
"111110001100000001110011000000000000",--8575
"001001111100000001001111111111111011",--8576
"001001111100000000111111111111111010",--8577
"001011111100000001101111111111111001",--8578
"001011111100000001011111111111111000",--8579
"001011111100000001001111111111110111",--8580
"001011111100000000111111111111110110",--8581
"101000000001111000000000100000000000",--8582
"101110001001111000000001100000000000",--8583
"101110001011111000000010000000000000",--8584
"101110001101111000000010100000000000",--8585
"001001111100000111111111111111110101",--8586
"101001111100010111100000000000001100",--8587
"000111000000000000000000011110001000",--8588
"101001111100000111100000000000001100",--8589
"001101111100000111111111111111110101",--8590
"010000000011000000000000000000001100",--8591
"001111111100000000111111111111110110",--8592
"001011000000000000110000000100101101",--8593
"001111111100000000111111111111110111",--8594
"001011000000000000110000000100101010",--8595
"001111111100000000111111111111111000",--8596
"001011000000000000110000000100101011",--8597
"001111111100000000111111111111111001",--8598
"001011000000000000110000000100101100",--8599
"001101111100000000011111111111111010",--8600
"001001000000000000010000000100101001",--8601
"001101111100000000011111111111111011",--8602
"001001000000000000010000000100101110",--8603
"101001000000000000010000000000000001",--8604
"001101111100000000101111111111111100",--8605
"001101111100000000110000000000000000",--8606
"001001111100000111111111111111111011",--8607
"101001111100010111100000000000000110",--8608
"000111000000000000000001011101010010",--8609
"101001111100000111100000000000000110",--8610
"001101111100000111111111111111111011",--8611
"001101111100000000011111111111111101",--8612
"001101000010000000100000000000000011",--8613
"010011000101000000000000001001010100",--8614
"001101000100000000100000000100110001",--8615
"001101111100000000110000000000000000",--8616
"101000000001111000000000100000000000",--8617
"001001111100000111111111111111111100",--8618
"101001111100010111100000000000000101",--8619
"000111000000000000000001011101010010",--8620
"101001111100000111100000000000000101",--8621
"101001000000000000010000000000000100",--8622
"001101111100000000101111111111111101",--8623
"001101111100000000110000000000000000",--8624
"101001111100010111100000000000000101",--8625
"000111000000000000000001110100010111",--8626
"101001111100000111100000000000000101",--8627
"001101111100000111111111111111111100",--8628
"000101000000000000000010001111111011",--8629
"001101001010000001010000000101101101",--8630
"001111000000000000110000000100010101",--8631
"001101001010000001100000000000000101",--8632
"001111001100000001000000000000000000",--8633
"111110000110010001000001100000000000",--8634
"001111000000000001000000000100010110",--8635
"001111001100000001010000000000000001",--8636
"111110001000010001010010000000000000",--8637
"001111000000000001010000000100010111",--8638
"001111001100000001100000000000000010",--8639
"111110001010010001100010100000000000",--8640
"001101001010000001100000000000000001",--8641
"011111001101000000010000000001010001",--8642
"001111000110000001100000000000000000",--8643
"010010001101000000000000000000011001",--8644
"001101001010000001100000000000000100",--8645
"001101001010000001110000000000000110",--8646
"011010001101000000000000000000000010",--8647
"101001000000000010000000000000000001",--8648
"000101000000000000000010000111001011",--8649
"101000000001111000000100000000000000",--8650
"001111001100000001100000000000000000",--8651
"011100001111000010000000000000000001",--8652
"101110001101111000000011000000000010",--8653
"111110001100010000110011000000000000",--8654
"001111000110000001110000000000000000",--8655
"111110001110011000000011100000000000",--8656
"111110001100001001110011000000000000",--8657
"001111000110000001110000000000000001",--8658
"111110001100001001110011100000000000",--8659
"111110001110000001000011100000000001",--8660
"001111001100000010000000000000000001",--8661
"010110010001000001110000000000000111",--8662
"001111000110000001110000000000000010",--8663
"111110001100001001110011100000000000",--8664
"111110001110000001010011100000000001",--8665
"001111001100000010000000000000000010",--8666
"010110010001000001110000000000000010",--8667
"001011000000000001100000000100101111",--8668
"000101000000000000000010001010100000",--8669
"001111000110000001100000000000000001",--8670
"010010001101000000000000000000011001",--8671
"001101001010000001100000000000000100",--8672
"001101001010000001110000000000000110",--8673
"011010001101000000000000000000000010",--8674
"101001000000000010000000000000000001",--8675
"000101000000000000000010000111100110",--8676
"101000000001111000000100000000000000",--8677
"001111001100000001100000000000000001",--8678
"011100001111000010000000000000000001",--8679
"101110001101111000000011000000000010",--8680
"111110001100010001000011000000000000",--8681
"001111000110000001110000000000000001",--8682
"111110001110011000000011100000000000",--8683
"111110001100001001110011000000000000",--8684
"001111000110000001110000000000000010",--8685
"111110001100001001110011100000000000",--8686
"111110001110000001010011100000000001",--8687
"001111001100000010000000000000000010",--8688
"010110010001000001110000000000000111",--8689
"001111000110000001110000000000000000",--8690
"111110001100001001110011100000000000",--8691
"111110001110000000110011100000000001",--8692
"001111001100000010000000000000000000",--8693
"010110010001000001110000000000000010",--8694
"001011000000000001100000000100101111",--8695
"000101000000000000000010001010100000",--8696
"001111000110000001100000000000000010",--8697
"010010001101000000000000001000000000",--8698
"001101001010000001100000000000000100",--8699
"001101001010000001010000000000000110",--8700
"011010001101000000000000000000000010",--8701
"101001000000000001110000000000000001",--8702
"000101000000000000000010001000000001",--8703
"101000000001111000000011100000000000",--8704
"001111001100000001100000000000000010",--8705
"011100001011000001110000000000000001",--8706
"101110001101111000000011000000000010",--8707
"111110001100010001010010100000000000",--8708
"001111000110000001100000000000000010",--8709
"111110001100011000000011000000000000",--8710
"111110001010001001100010100000000000",--8711
"001111000110000001100000000000000000",--8712
"111110001010001001100011000000000000",--8713
"111110001100000000110001100000000001",--8714
"001111001100000001100000000000000000",--8715
"010110001101000000110000000111101110",--8716
"001111000110000000110000000000000001",--8717
"111110001010001000110001100000000000",--8718
"111110000110000001000001100000000001",--8719
"001111001100000001000000000000000001",--8720
"010110001001000000110000000111101001",--8721
"001011000000000001010000000100101111",--8722
"000101000000000000000010001010100000",--8723
"011111001101000000100000000000011001",--8724
"001101001010000001010000000000000100",--8725
"001111000110000001100000000000000000",--8726
"001111001010000001110000000000000000",--8727
"111110001100001001110011000000000000",--8728
"001111000110000001110000000000000001",--8729
"001111001010000010000000000000000001",--8730
"111110001110001010000011100000000000",--8731
"111110001100000001110011000000000000",--8732
"001111000110000001110000000000000010",--8733
"001111001010000010000000000000000010",--8734
"111110001110001010000011100000000000",--8735
"111110001100000001110011000000000000",--8736
"010110001101000000000000000111011001",--8737
"001111001010000001110000000000000000",--8738
"111110001110001000110001100000000000",--8739
"001111001010000001110000000000000001",--8740
"111110001110001001000010000000000000",--8741
"111110000110000001000001100000000000",--8742
"001111001010000001000000000000000010",--8743
"111110001000001001010010000000000000",--8744
"111110000110000001000001100000000010",--8745
"111110001100011000000010000000000000",--8746
"111110000110001001000001100000000000",--8747
"001011000000000000110000000100101111",--8748
"000101000000000000000010001010100000",--8749
"001111000110000001100000000000000000",--8750
"001111000110000001110000000000000001",--8751
"001111000110000010000000000000000010",--8752
"111110001100001001100100100000000000",--8753
"001101001010000001110000000000000100",--8754
"001111001110000010100000000000000000",--8755
"111110010010001010100100100000000000",--8756
"111110001110001001110101000000000000",--8757
"001111001110000010110000000000000001",--8758
"111110010100001010110101000000000000",--8759
"111110010010000010100100100000000000",--8760
"111110010000001010000101000000000000",--8761
"001111001110000010110000000000000010",--8762
"111110010100001010110101000000000000",--8763
"111110010010000010100100100000000000",--8764
"001101001010000010000000000000000011",--8765
"011100010001000000000000000000000011",--8766
"101110010011111000000011000000000000",--8767
"011110010011000000000000000000001111",--8768
"000101000000000000000010001111111011",--8769
"111110001110001010000101000000000000",--8770
"001101001010000010010000000000001001",--8771
"001111010010000010110000000000000000",--8772
"111110010100001010110101000000000000",--8773
"111110010010000010100100100000000000",--8774
"111110010000001001100100000000000000",--8775
"001111010010000010100000000000000001",--8776
"111110010000001010100100000000000000",--8777
"111110010010000010000100000000000000",--8778
"111110001100001001110011000000000000",--8779
"001111010010000001110000000000000010",--8780
"111110001100001001110011000000000000",--8781
"111110010000000001100011000000000000",--8782
"010010001101000000000000000110101011",--8783
"001111000110000001110000000000000000",--8784
"001111000110000010000000000000000001",--8785
"001111000110000010010000000000000010",--8786
"111110001110001000110101000000000000",--8787
"001111001110000010110000000000000000",--8788
"111110010100001010110101000000000000",--8789
"111110010000001001000101100000000000",--8790
"001111001110000011000000000000000001",--8791
"111110010110001011000101100000000000",--8792
"111110010100000010110101000000000000",--8793
"111110010010001001010101100000000000",--8794
"001111001110000011000000000000000010",--8795
"111110010110001011000101100000000000",--8796
"111110010100000010110101000000000000",--8797
"011100010001000000000000000000000010",--8798
"101110010101111000000011100000000000",--8799
"000101000000000000000010001001110110",--8800
"111110010010001001000101100000000000",--8801
"111110010000001001010110000000000000",--8802
"111110010110000011000101100000000000",--8803
"001101001010000010010000000000001001",--8804
"001111010010000011000000000000000000",--8805
"111110010110001011000101100000000000",--8806
"111110001110001001010110000000000000",--8807
"111110010010001000110100100000000000",--8808
"111110011000000010010100100000000000",--8809
"001111010010000011000000000000000001",--8810
"111110010010001011000100100000000000",--8811
"111110010110000010010100100000000000",--8812
"111110001110001001000011100000000000",--8813
"111110010000001000110100000000000000",--8814
"111110001110000010000011100000000000",--8815
"001111010010000010000000000000000010",--8816
"111110001110001010000011100000000000",--8817
"111110010010000001110011100000000000",--8818
"101111000001110010000011111100000000",--8819
"111110001110001010000011100000000000",--8820
"111110010100000001110011100000000000",--8821
"111110000110001000110100000000000000",--8822
"001111001110000010010000000000000000",--8823
"111110010000001010010100000000000000",--8824
"111110001000001001000100100000000000",--8825
"001111001110000010100000000000000001",--8826
"111110010010001010100100100000000000",--8827
"111110010000000010010100000000000000",--8828
"111110001010001001010100100000000000",--8829
"001111001110000010100000000000000010",--8830
"111110010010001010100100100000000000",--8831
"111110010000000010010100000000000000",--8832
"011100010001000000000000000000000011",--8833
"101110010001111000000001100000000000",--8834
"011111001101000000110000000000010000",--8835
"000101000000000000000010001010010011",--8836
"111110001000001001010100100000000000",--8837
"001101001010000001110000000000001001",--8838
"001111001110000010100000000000000000",--8839
"111110010010001010100100100000000000",--8840
"111110010000000010010100000000000000",--8841
"111110001010001000110010100000000000",--8842
"001111001110000010010000000000000001",--8843
"111110001010001010010010100000000000",--8844
"111110010000000001010010100000000000",--8845
"111110000110001001000001100000000000",--8846
"001111001110000001000000000000000010",--8847
"111110000110001001000001100000000000",--8848
"111110001010000000110001100000000000",--8849
"011111001101000000110000000000000001",--8850
"111110000110010000010001100000000000",--8851
"111110001110001001110010000000000000",--8852
"111110001100001000110001100000000000",--8853
"111110001000010000110001100000000000",--8854
"010110000111000000000000000101100011",--8855
"111110000110100000000001100000000000",--8856
"001101001010000001010000000000000110",--8857
"011100001011000000000000000000000001",--8858
"101110000111111000000001100000000010",--8859
"111110000110010001110001100000000000",--8860
"111110001100011000000010000000000000",--8861
"111110000110001001000001100000000000",--8862
"001011000000000000110000000100101111",--8863
"001111000000000000110000000100101111",--8864
"001111000000000001000000000100101101",--8865
"010110001001000000110000000101011000",--8866
"001101001000000001010000000000000001",--8867
"010011001011000000000000000101010110",--8868
"001101001010000000100000000100110001",--8869
"001001111100000001001111111111111101",--8870
"101000000001111000000000100000000000",--8871
"001001111100000111111111111111111100",--8872
"101001111100010111100000000000000101",--8873
"000111000000000000000001011101010010",--8874
"101001111100000111100000000000000101",--8875
"001101111100000111111111111111111100",--8876
"001101111100000000011111111111111101",--8877
"001101000010000000100000000000000010",--8878
"010011000101000000000000000101001011",--8879
"001101000100000000100000000100110001",--8880
"001101000100000000110000000000000000",--8881
"010011000111000000000000000100110111",--8882
"001101000110000001000000000101101101",--8883
"001111000000000000110000000100010101",--8884
"001101001000000001010000000000000101",--8885
"001111001010000001000000000000000000",--8886
"111110000110010001000001100000000000",--8887
"001111000000000001000000000100010110",--8888
"001111001010000001010000000000000001",--8889
"111110001000010001010010000000000000",--8890
"001111000000000001010000000100010111",--8891
"001111001010000001100000000000000010",--8892
"111110001010010001100010100000000000",--8893
"001101001000000001010000000000000001",--8894
"011111001011000000010000000001010101",--8895
"001101111100000001010000000000000000",--8896
"001111001010000001100000000000000000",--8897
"010010001101000000000000000000011010",--8898
"001101001000000001100000000000000100",--8899
"001101001000000001110000000000000110",--8900
"011010001101000000000000000000000010",--8901
"101001000000000010000000000000000001",--8902
"000101000000000000000010001011001001",--8903
"101000000001111000000100000000000000",--8904
"001111001100000001100000000000000000",--8905
"011100001111000010000000000000000001",--8906
"101110001101111000000011000000000010",--8907
"111110001100010000110011000000000000",--8908
"001111001010000001110000000000000000",--8909
"111110001110011000000011100000000000",--8910
"111110001100001001110011000000000000",--8911
"001111001010000001110000000000000001",--8912
"111110001100001001110011100000000000",--8913
"111110001110000001000011100000000001",--8914
"001111001100000010000000000000000001",--8915
"010110010001000001110000000000001000",--8916
"001111001010000001110000000000000010",--8917
"111110001100001001110011100000000000",--8918
"111110001110000001010011100000000001",--8919
"001111001100000010000000000000000010",--8920
"010110010001000001110000000000000011",--8921
"001011000000000001100000000100101111",--8922
"101001000000000001000000000000000001",--8923
"000101000000000000000010001110110001",--8924
"001111001010000001100000000000000001",--8925
"010010001101000000000000000000011010",--8926
"001101001000000001100000000000000100",--8927
"001101001000000001110000000000000110",--8928
"011010001101000000000000000000000010",--8929
"101001000000000010000000000000000001",--8930
"000101000000000000000010001011100101",--8931
"101000000001111000000100000000000000",--8932
"001111001100000001100000000000000001",--8933
"011100001111000010000000000000000001",--8934
"101110001101111000000011000000000010",--8935
"111110001100010001000011000000000000",--8936
"001111001010000001110000000000000001",--8937
"111110001110011000000011100000000000",--8938
"111110001100001001110011000000000000",--8939
"001111001010000001110000000000000010",--8940
"111110001100001001110011100000000000",--8941
"111110001110000001010011100000000001",--8942
"001111001100000010000000000000000010",--8943
"010110010001000001110000000000001000",--8944
"001111001010000001110000000000000000",--8945
"111110001100001001110011100000000000",--8946
"111110001110000000110011100000000001",--8947
"001111001100000010000000000000000000",--8948
"010110010001000001110000000000000011",--8949
"001011000000000001100000000100101111",--8950
"101001000000000001000000000000000010",--8951
"000101000000000000000010001110110001",--8952
"001111001010000001100000000000000010",--8953
"010010001101000000000000000010101011",--8954
"001101001000000001100000000000000100",--8955
"001101001000000001000000000000000110",--8956
"011010001101000000000000000000000010",--8957
"101001000000000001110000000000000001",--8958
"000101000000000000000010001100000001",--8959
"101000000001111000000011100000000000",--8960
"001111001100000001100000000000000010",--8961
"011100001001000001110000000000000001",--8962
"101110001101111000000011000000000010",--8963
"111110001100010001010010100000000000",--8964
"001111001010000001100000000000000010",--8965
"111110001100011000000011000000000000",--8966
"111110001010001001100010100000000000",--8967
"001111001010000001100000000000000000",--8968
"111110001010001001100011000000000000",--8969
"111110001100000000110001100000000001",--8970
"001111001100000001100000000000000000",--8971
"010110001101000000110000000010011001",--8972
"001111001010000000110000000000000001",--8973
"111110001010001000110001100000000000",--8974
"111110000110000001000001100000000001",--8975
"001111001100000001000000000000000001",--8976
"010110001001000000110000000010010100",--8977
"001011000000000001010000000100101111",--8978
"101001000000000001000000000000000011",--8979
"000101000000000000000010001110110001",--8980
"011111001011000000100000000000011011",--8981
"001101001000000001000000000000000100",--8982
"001101111100000001010000000000000000",--8983
"001111001010000001100000000000000000",--8984
"001111001000000001110000000000000000",--8985
"111110001100001001110011000000000000",--8986
"001111001010000001110000000000000001",--8987
"001111001000000010000000000000000001",--8988
"111110001110001010000011100000000000",--8989
"111110001100000001110011000000000000",--8990
"001111001010000001110000000000000010",--8991
"001111001000000010000000000000000010",--8992
"111110001110001010000011100000000000",--8993
"111110001100000001110011000000000000",--8994
"010110001101000000000000000010000010",--8995
"001111001000000001110000000000000000",--8996
"111110001110001000110001100000000000",--8997
"001111001000000001110000000000000001",--8998
"111110001110001001000010000000000000",--8999
"111110000110000001000001100000000000",--9000
"001111001000000001000000000000000010",--9001
"111110001000001001010010000000000000",--9002
"111110000110000001000001100000000010",--9003
"111110001100011000000010000000000000",--9004
"111110000110001001000001100000000000",--9005
"001011000000000000110000000100101111",--9006
"101001000000000001000000000000000001",--9007
"000101000000000000000010001110110001",--9008
"001101111100000001100000000000000000",--9009
"001111001100000001100000000000000000",--9010
"001111001100000001110000000000000001",--9011
"001111001100000010000000000000000010",--9012
"111110001100001001100100100000000000",--9013
"001101001000000001110000000000000100",--9014
"001111001110000010100000000000000000",--9015
"111110010010001010100100100000000000",--9016
"111110001110001001110101000000000000",--9017
"001111001110000010110000000000000001",--9018
"111110010100001010110101000000000000",--9019
"111110010010000010100100100000000000",--9020
"111110010000001010000101000000000000",--9021
"001111001110000010110000000000000010",--9022
"111110010100001010110101000000000000",--9023
"111110010010000010100100100000000000",--9024
"001101001000000010000000000000000011",--9025
"011100010001000000000000000000000011",--9026
"101110010011111000000011000000000000",--9027
"011110010011000000000000000000001111",--9028
"000101000000000000000010001110100110",--9029
"111110001110001010000101000000000000",--9030
"001101001000000010010000000000001001",--9031
"001111010010000010110000000000000000",--9032
"111110010100001010110101000000000000",--9033
"111110010010000010100100100000000000",--9034
"111110010000001001100100000000000000",--9035
"001111010010000010100000000000000001",--9036
"111110010000001010100100000000000000",--9037
"111110010010000010000100000000000000",--9038
"111110001100001001110011000000000000",--9039
"001111010010000001110000000000000010",--9040
"111110001100001001110011000000000000",--9041
"111110010000000001100011000000000000",--9042
"010010001101000000000000000001010010",--9043
"001111001100000001110000000000000000",--9044
"001111001100000010000000000000000001",--9045
"001111001100000010010000000000000010",--9046
"111110001110001000110101000000000000",--9047
"001111001110000010110000000000000000",--9048
"111110010100001010110101000000000000",--9049
"111110010000001001000101100000000000",--9050
"001111001110000011000000000000000001",--9051
"111110010110001011000101100000000000",--9052
"111110010100000010110101000000000000",--9053
"111110010010001001010101100000000000",--9054
"001111001110000011000000000000000010",--9055
"111110010110001011000101100000000000",--9056
"111110010100000010110101000000000000",--9057
"011100010001000000000000000000000010",--9058
"101110010101111000000011100000000000",--9059
"000101000000000000000010001101111010",--9060
"111110010010001001000101100000000000",--9061
"111110010000001001010110000000000000",--9062
"111110010110000011000101100000000000",--9063
"001101001000000010010000000000001001",--9064
"001111010010000011000000000000000000",--9065
"111110010110001011000101100000000000",--9066
"111110001110001001010110000000000000",--9067
"111110010010001000110100100000000000",--9068
"111110011000000010010100100000000000",--9069
"001111010010000011000000000000000001",--9070
"111110010010001011000100100000000000",--9071
"111110010110000010010100100000000000",--9072
"111110001110001001000011100000000000",--9073
"111110010000001000110100000000000000",--9074
"111110001110000010000011100000000000",--9075
"001111010010000010000000000000000010",--9076
"111110001110001010000011100000000000",--9077
"111110010010000001110011100000000000",--9078
"101111000001110010000011111100000000",--9079
"111110001110001010000011100000000000",--9080
"111110010100000001110011100000000000",--9081
"111110000110001000110100000000000000",--9082
"001111001110000010010000000000000000",--9083
"111110010000001010010100000000000000",--9084
"111110001000001001000100100000000000",--9085
"001111001110000010100000000000000001",--9086
"111110010010001010100100100000000000",--9087
"111110010000000010010100000000000000",--9088
"111110001010001001010100100000000000",--9089
"001111001110000010100000000000000010",--9090
"111110010010001010100100100000000000",--9091
"111110010000000010010100000000000000",--9092
"011100010001000000000000000000000011",--9093
"101110010001111000000001100000000000",--9094
"011111001011000000110000000000010000",--9095
"000101000000000000000010001110010111",--9096
"111110001000001001010100100000000000",--9097
"001101001000000001110000000000001001",--9098
"001111001110000010100000000000000000",--9099
"111110010010001010100100100000000000",--9100
"111110010000000010010100000000000000",--9101
"111110001010001000110010100000000000",--9102
"001111001110000010010000000000000001",--9103
"111110001010001010010010100000000000",--9104
"111110010000000001010010100000000000",--9105
"111110000110001001000001100000000000",--9106
"001111001110000001000000000000000010",--9107
"111110000110001001000001100000000000",--9108
"111110001010000000110001100000000000",--9109
"011111001011000000110000000000000001",--9110
"111110000110010000010001100000000000",--9111
"111110001110001001110010000000000000",--9112
"111110001100001000110001100000000000",--9113
"111110001000010000110001100000000000",--9114
"010110000111000000000000000000001010",--9115
"111110000110100000000001100000000000",--9116
"001101001000000001000000000000000110",--9117
"011100001001000000000000000000000001",--9118
"101110000111111000000001100000000010",--9119
"111110000110010001110001100000000000",--9120
"111110001100011000000010000000000000",--9121
"111110000110001001000001100000000000",--9122
"001011000000000000110000000100101111",--9123
"101001000000000001000000000000000001",--9124
"000101000000000000000010001110110001",--9125
"001101000110000000110000000101101101",--9126
"001101000110000000110000000000000110",--9127
"010000000111000000000000000001000001",--9128
"001101111100000000110000000000000000",--9129
"101001000000000000010000000000000001",--9130
"001001111100000111111111111111111100",--9131
"101001111100010111100000000000000101",--9132
"000111000000000000000001011101010010",--9133
"101001111100000111100000000000000101",--9134
"001101111100000111111111111111111100",--9135
"000101000000000000000010001111101010",--9136
"001111000000000000110000000100101111",--9137
"001001111100000000101111111111111100",--9138
"010110000111000000000000000000101110",--9139
"001111000000000001000000000100101101",--9140
"010110001001000000110000000000101100",--9141
"101111001001110001000011110000100011",--9142
"101111001001100001001101011100001010",--9143
"111110000110000001000001100000000000",--9144
"001101111100000001010000000000000000",--9145
"001111001010000001000000000000000000",--9146
"111110001000001000110010000000000000",--9147
"001111000000000001010000000100010101",--9148
"111110001000000001010010000000000000",--9149
"001111001010000001010000000000000001",--9150
"111110001010001000110010100000000000",--9151
"001111000000000001100000000100010110",--9152
"111110001010000001100010100000000000",--9153
"001111001010000001100000000000000010",--9154
"111110001100001000110011000000000000",--9155
"001111000000000001110000000100010111",--9156
"111110001100000001110011000000000000",--9157
"001001111100000001001111111111111011",--9158
"001001111100000000111111111111111010",--9159
"001011111100000001101111111111111001",--9160
"001011111100000001011111111111111000",--9161
"001011111100000001001111111111110111",--9162
"001011111100000000111111111111110110",--9163
"101000000001111000000000100000000000",--9164
"101110001001111000000001100000000000",--9165
"101110001011111000000010000000000000",--9166
"101110001101111000000010100000000000",--9167
"001001111100000111111111111111110101",--9168
"101001111100010111100000000000001100",--9169
"000111000000000000000000011110001000",--9170
"101001111100000111100000000000001100",--9171
"001101111100000111111111111111110101",--9172
"010000000011000000000000000000001100",--9173
"001111111100000000111111111111110110",--9174
"001011000000000000110000000100101101",--9175
"001111111100000000111111111111110111",--9176
"001011000000000000110000000100101010",--9177
"001111111100000000111111111111111000",--9178
"001011000000000000110000000100101011",--9179
"001111111100000000111111111111111001",--9180
"001011000000000000110000000100101100",--9181
"001101111100000000011111111111111010",--9182
"001001000000000000010000000100101001",--9183
"001101111100000000011111111111111011",--9184
"001001000000000000010000000100101110",--9185
"101001000000000000010000000000000001",--9186
"001101111100000000101111111111111100",--9187
"001101111100000000110000000000000000",--9188
"001001111100000111111111111111111011",--9189
"101001111100010111100000000000000110",--9190
"000111000000000000000001011101010010",--9191
"101001111100000111100000000000000110",--9192
"001101111100000111111111111111111011",--9193
"001101111100000000011111111111111101",--9194
"001101000010000000100000000000000011",--9195
"010011000101000000000000000000001110",--9196
"001101000100000000100000000100110001",--9197
"001101111100000000110000000000000000",--9198
"101000000001111000000000100000000000",--9199
"001001111100000111111111111111111100",--9200
"101001111100010111100000000000000101",--9201
"000111000000000000000001011101010010",--9202
"101001111100000111100000000000000101",--9203
"101001000000000000010000000000000100",--9204
"001101111100000000101111111111111101",--9205
"001101111100000000110000000000000000",--9206
"101001111100010111100000000000000101",--9207
"000111000000000000000001110100010111",--9208
"101001111100000111100000000000000101",--9209
"001101111100000111111111111111111100",--9210
"001101111100000000011111111111111110",--9211
"101001000010000000010000000000000001",--9212
"001101111100000000111111111111111111",--9213
"001100000110000000010001000000000000",--9214
"001101000100000001000000000000000000",--9215
"010011001000000000001111100000000000",--9216
"001001111100000000011111111111111101",--9217
"011111001001011000110000000101010001",--9218
"001101000100000001000000000000000001",--9219
"010011001001000000000000001110001111",--9220
"001101001000000001000000000100110001",--9221
"001101001000000001010000000000000000",--9222
"001001111100000000101111111111111100",--9223
"010011001011000000000000000100111001",--9224
"001101001010000001100000000101101101",--9225
"001111000000000000110000000100010101",--9226
"001101001100000001110000000000000101",--9227
"001111001110000001000000000000000000",--9228
"111110000110010001000001100000000000",--9229
"001111000000000001000000000100010110",--9230
"001111001110000001010000000000000001",--9231
"111110001000010001010010000000000000",--9232
"001111000000000001010000000100010111",--9233
"001111001110000001100000000000000010",--9234
"111110001010010001100010100000000000",--9235
"001101001100000001110000000000000001",--9236
"011111001111000000010000000001010101",--9237
"001101111100000001110000000000000000",--9238
"001111001110000001100000000000000000",--9239
"010010001101000000000000000000011010",--9240
"001101001100000010000000000000000100",--9241
"001101001100000010010000000000000110",--9242
"011010001101000000000000000000000010",--9243
"101001000000000010100000000000000001",--9244
"000101000000000000000010010000011111",--9245
"101000000001111000000101000000000000",--9246
"001111010000000001100000000000000000",--9247
"011100010011000010100000000000000001",--9248
"101110001101111000000011000000000010",--9249
"111110001100010000110011000000000000",--9250
"001111001110000001110000000000000000",--9251
"111110001110011000000011100000000000",--9252
"111110001100001001110011000000000000",--9253
"001111001110000001110000000000000001",--9254
"111110001100001001110011100000000000",--9255
"111110001110000001000011100000000001",--9256
"001111010000000010000000000000000001",--9257
"010110010001000001110000000000001000",--9258
"001111001110000001110000000000000010",--9259
"111110001100001001110011100000000000",--9260
"111110001110000001010011100000000001",--9261
"001111010000000010000000000000000010",--9262
"010110010001000001110000000000000011",--9263
"001011000000000001100000000100101111",--9264
"101001000000000001100000000000000001",--9265
"000101000000000000000010010100001000",--9266
"001111001110000001100000000000000001",--9267
"010010001101000000000000000000011010",--9268
"001101001100000010000000000000000100",--9269
"001101001100000010010000000000000110",--9270
"011010001101000000000000000000000010",--9271
"101001000000000010100000000000000001",--9272
"000101000000000000000010010000111011",--9273
"101000000001111000000101000000000000",--9274
"001111010000000001100000000000000001",--9275
"011100010011000010100000000000000001",--9276
"101110001101111000000011000000000010",--9277
"111110001100010001000011000000000000",--9278
"001111001110000001110000000000000001",--9279
"111110001110011000000011100000000000",--9280
"111110001100001001110011000000000000",--9281
"001111001110000001110000000000000010",--9282
"111110001100001001110011100000000000",--9283
"111110001110000001010011100000000001",--9284
"001111010000000010000000000000000010",--9285
"010110010001000001110000000000001000",--9286
"001111001110000001110000000000000000",--9287
"111110001100001001110011100000000000",--9288
"111110001110000000110011100000000001",--9289
"001111010000000010000000000000000000",--9290
"010110010001000001110000000000000011",--9291
"001011000000000001100000000100101111",--9292
"101001000000000001100000000000000010",--9293
"000101000000000000000010010100001000",--9294
"001111001110000001100000000000000010",--9295
"010010001101000000000000000010101011",--9296
"001101001100000010000000000000000100",--9297
"001101001100000001100000000000000110",--9298
"011010001101000000000000000000000010",--9299
"101001000000000010010000000000000001",--9300
"000101000000000000000010010001010111",--9301
"101000000001111000000100100000000000",--9302
"001111010000000001100000000000000010",--9303
"011100001101000010010000000000000001",--9304
"101110001101111000000011000000000010",--9305
"111110001100010001010010100000000000",--9306
"001111001110000001100000000000000010",--9307
"111110001100011000000011000000000000",--9308
"111110001010001001100010100000000000",--9309
"001111001110000001100000000000000000",--9310
"111110001010001001100011000000000000",--9311
"111110001100000000110001100000000001",--9312
"001111010000000001100000000000000000",--9313
"010110001101000000110000000010011001",--9314
"001111001110000000110000000000000001",--9315
"111110001010001000110001100000000000",--9316
"111110000110000001000001100000000001",--9317
"001111010000000001000000000000000001",--9318
"010110001001000000110000000010010100",--9319
"001011000000000001010000000100101111",--9320
"101001000000000001100000000000000011",--9321
"000101000000000000000010010100001000",--9322
"011111001111000000100000000000011011",--9323
"001101001100000001100000000000000100",--9324
"001101111100000001110000000000000000",--9325
"001111001110000001100000000000000000",--9326
"001111001100000001110000000000000000",--9327
"111110001100001001110011000000000000",--9328
"001111001110000001110000000000000001",--9329
"001111001100000010000000000000000001",--9330
"111110001110001010000011100000000000",--9331
"111110001100000001110011000000000000",--9332
"001111001110000001110000000000000010",--9333
"001111001100000010000000000000000010",--9334
"111110001110001010000011100000000000",--9335
"111110001100000001110011000000000000",--9336
"010110001101000000000000000010000010",--9337
"001111001100000001110000000000000000",--9338
"111110001110001000110001100000000000",--9339
"001111001100000001110000000000000001",--9340
"111110001110001001000010000000000000",--9341
"111110000110000001000001100000000000",--9342
"001111001100000001000000000000000010",--9343
"111110001000001001010010000000000000",--9344
"111110000110000001000001100000000010",--9345
"111110001100011000000010000000000000",--9346
"111110000110001001000001100000000000",--9347
"001011000000000000110000000100101111",--9348
"101001000000000001100000000000000001",--9349
"000101000000000000000010010100001000",--9350
"001101111100000010000000000000000000",--9351
"001111010000000001100000000000000000",--9352
"001111010000000001110000000000000001",--9353
"001111010000000010000000000000000010",--9354
"111110001100001001100100100000000000",--9355
"001101001100000010010000000000000100",--9356
"001111010010000010100000000000000000",--9357
"111110010010001010100100100000000000",--9358
"111110001110001001110101000000000000",--9359
"001111010010000010110000000000000001",--9360
"111110010100001010110101000000000000",--9361
"111110010010000010100100100000000000",--9362
"111110010000001010000101000000000000",--9363
"001111010010000010110000000000000010",--9364
"111110010100001010110101000000000000",--9365
"111110010010000010100100100000000000",--9366
"001101001100000010100000000000000011",--9367
"011100010101000000000000000000000011",--9368
"101110010011111000000011000000000000",--9369
"011110010011000000000000000000001111",--9370
"000101000000000000000010010011111100",--9371
"111110001110001010000101000000000000",--9372
"001101001100000010110000000000001001",--9373
"001111010110000010110000000000000000",--9374
"111110010100001010110101000000000000",--9375
"111110010010000010100100100000000000",--9376
"111110010000001001100100000000000000",--9377
"001111010110000010100000000000000001",--9378
"111110010000001010100100000000000000",--9379
"111110010010000010000100000000000000",--9380
"111110001100001001110011000000000000",--9381
"001111010110000001110000000000000010",--9382
"111110001100001001110011000000000000",--9383
"111110010000000001100011000000000000",--9384
"010010001101000000000000000001010010",--9385
"001111010000000001110000000000000000",--9386
"001111010000000010000000000000000001",--9387
"001111010000000010010000000000000010",--9388
"111110001110001000110101000000000000",--9389
"001111010010000010110000000000000000",--9390
"111110010100001010110101000000000000",--9391
"111110010000001001000101100000000000",--9392
"001111010010000011000000000000000001",--9393
"111110010110001011000101100000000000",--9394
"111110010100000010110101000000000000",--9395
"111110010010001001010101100000000000",--9396
"001111010010000011000000000000000010",--9397
"111110010110001011000101100000000000",--9398
"111110010100000010110101000000000000",--9399
"011100010101000000000000000000000010",--9400
"101110010101111000000011100000000000",--9401
"000101000000000000000010010011010000",--9402
"111110010010001001000101100000000000",--9403
"111110010000001001010110000000000000",--9404
"111110010110000011000101100000000000",--9405
"001101001100000010110000000000001001",--9406
"001111010110000011000000000000000000",--9407
"111110010110001011000101100000000000",--9408
"111110001110001001010110000000000000",--9409
"111110010010001000110100100000000000",--9410
"111110011000000010010100100000000000",--9411
"001111010110000011000000000000000001",--9412
"111110010010001011000100100000000000",--9413
"111110010110000010010100100000000000",--9414
"111110001110001001000011100000000000",--9415
"111110010000001000110100000000000000",--9416
"111110001110000010000011100000000000",--9417
"001111010110000010000000000000000010",--9418
"111110001110001010000011100000000000",--9419
"111110010010000001110011100000000000",--9420
"101111000001110010000011111100000000",--9421
"111110001110001010000011100000000000",--9422
"111110010100000001110011100000000000",--9423
"111110000110001000110100000000000000",--9424
"001111010010000010010000000000000000",--9425
"111110010000001010010100000000000000",--9426
"111110001000001001000100100000000000",--9427
"001111010010000010100000000000000001",--9428
"111110010010001010100100100000000000",--9429
"111110010000000010010100000000000000",--9430
"111110001010001001010100100000000000",--9431
"001111010010000010100000000000000010",--9432
"111110010010001010100100100000000000",--9433
"111110010000000010010100000000000000",--9434
"011100010101000000000000000000000011",--9435
"101110010001111000000001100000000000",--9436
"011111001111000000110000000000010000",--9437
"000101000000000000000010010011101101",--9438
"111110001000001001010100100000000000",--9439
"001101001100000010010000000000001001",--9440
"001111010010000010100000000000000000",--9441
"111110010010001010100100100000000000",--9442
"111110010000000010010100000000000000",--9443
"111110001010001000110010100000000000",--9444
"001111010010000010010000000000000001",--9445
"111110001010001010010010100000000000",--9446
"111110010000000001010010100000000000",--9447
"111110000110001001000001100000000000",--9448
"001111010010000001000000000000000010",--9449
"111110000110001001000001100000000000",--9450
"111110001010000000110001100000000000",--9451
"011111001111000000110000000000000001",--9452
"111110000110010000010001100000000000",--9453
"111110001110001001110010000000000000",--9454
"111110001100001000110001100000000000",--9455
"111110001000010000110001100000000000",--9456
"010110000111000000000000000000001010",--9457
"111110000110100000000001100000000000",--9458
"001101001100000001100000000000000110",--9459
"011100001101000000000000000000000001",--9460
"101110000111111000000001100000000010",--9461
"111110000110010001110001100000000000",--9462
"111110001100011000000010000000000000",--9463
"111110000110001001000001100000000000",--9464
"001011000000000000110000000100101111",--9465
"101001000000000001100000000000000001",--9466
"000101000000000000000010010100001000",--9467
"001101001010000001010000000101101101",--9468
"001101001010000001010000000000000110",--9469
"010000001011000000000000000001000011",--9470
"001101111100000000110000000000000000",--9471
"101000001001111000000001000000000000",--9472
"101001000000000000010000000000000001",--9473
"001001111100000111111111111111111011",--9474
"101001111100010111100000000000000110",--9475
"000111000000000000000001011101010010",--9476
"101001111100000111100000000000000110",--9477
"001101111100000111111111111111111011",--9478
"000101000000000000000010010101000010",--9479
"001111000000000000110000000100101111",--9480
"001001111100000001001111111111111011",--9481
"010110000111000000000000000000101111",--9482
"001111000000000001000000000100101101",--9483
"010110001001000000110000000000101101",--9484
"101111001001110001000011110000100011",--9485
"101111001001100001001101011100001010",--9486
"111110000110000001000001100000000000",--9487
"001101111100000001110000000000000000",--9488
"001111001110000001000000000000000000",--9489
"111110001000001000110010000000000000",--9490
"001111000000000001010000000100010101",--9491
"111110001000000001010010000000000000",--9492
"001111001110000001010000000000000001",--9493
"111110001010001000110010100000000000",--9494
"001111000000000001100000000100010110",--9495
"111110001010000001100010100000000000",--9496
"001111001110000001100000000000000010",--9497
"111110001100001000110011000000000000",--9498
"001111000000000001110000000100010111",--9499
"111110001100000001110011000000000000",--9500
"001001111100000001101111111111111010",--9501
"001001111100000001011111111111111001",--9502
"001011111100000001101111111111111000",--9503
"001011111100000001011111111111110111",--9504
"001011111100000001001111111111110110",--9505
"001011111100000000111111111111110101",--9506
"101000001001111000000001000000000000",--9507
"101000000001111000000000100000000000",--9508
"101110001001111000000001100000000000",--9509
"101110001011111000000010000000000000",--9510
"101110001101111000000010100000000000",--9511
"001001111100000111111111111111110100",--9512
"101001111100010111100000000000001101",--9513
"000111000000000000000000011110001000",--9514
"101001111100000111100000000000001101",--9515
"001101111100000111111111111111110100",--9516
"010000000011000000000000000000001100",--9517
"001111111100000000111111111111110101",--9518
"001011000000000000110000000100101101",--9519
"001111111100000000111111111111110110",--9520
"001011000000000000110000000100101010",--9521
"001111111100000000111111111111110111",--9522
"001011000000000000110000000100101011",--9523
"001111111100000000111111111111111000",--9524
"001011000000000000110000000100101100",--9525
"001101111100000000011111111111111001",--9526
"001001000000000000010000000100101001",--9527
"001101111100000000011111111111111010",--9528
"001001000000000000010000000100101110",--9529
"101001000000000000010000000000000001",--9530
"001101111100000000101111111111111011",--9531
"001101111100000000110000000000000000",--9532
"001001111100000111111111111111111010",--9533
"101001111100010111100000000000000111",--9534
"000111000000000000000001011101010010",--9535
"101001111100000111100000000000000111",--9536
"001101111100000111111111111111111010",--9537
"001101111100000000011111111111111100",--9538
"001101000010000000100000000000000010",--9539
"010011000101000000000000001001001111",--9540
"001101000100000000100000000100110001",--9541
"001101111100000000110000000000000000",--9542
"101000000001111000000000100000000000",--9543
"001001111100000111111111111111111011",--9544
"101001111100010111100000000000000110",--9545
"000111000000000000000001011101010010",--9546
"101001111100000111100000000000000110",--9547
"101001000000000000010000000000000011",--9548
"001101111100000000101111111111111100",--9549
"001101111100000000110000000000000000",--9550
"101001111100010111100000000000000110",--9551
"000111000000000000000001110100010111",--9552
"101001111100000111100000000000000110",--9553
"001101111100000111111111111111111011",--9554
"000101000000000000000010011110010100",--9555
"001101001000000001000000000101101101",--9556
"001111000000000000110000000100010101",--9557
"001101001000000001010000000000000101",--9558
"001111001010000001000000000000000000",--9559
"111110000110010001000001100000000000",--9560
"001111000000000001000000000100010110",--9561
"001111001010000001010000000000000001",--9562
"111110001000010001010010000000000000",--9563
"001111000000000001010000000100010111",--9564
"001111001010000001100000000000000010",--9565
"111110001010010001100010100000000000",--9566
"001101001000000001010000000000000001",--9567
"011111001011000000010000000001010010",--9568
"001101111100000001010000000000000000",--9569
"001111001010000001100000000000000000",--9570
"010010001101000000000000000000011001",--9571
"001101001000000001100000000000000100",--9572
"001101001000000001110000000000000110",--9573
"011010001101000000000000000000000010",--9574
"101001000000000010000000000000000001",--9575
"000101000000000000000010010101101010",--9576
"101000000001111000000100000000000000",--9577
"001111001100000001100000000000000000",--9578
"011100001111000010000000000000000001",--9579
"101110001101111000000011000000000010",--9580
"111110001100010000110011000000000000",--9581
"001111001010000001110000000000000000",--9582
"111110001110011000000011100000000000",--9583
"111110001100001001110011000000000000",--9584
"001111001010000001110000000000000001",--9585
"111110001100001001110011100000000000",--9586
"111110001110000001000011100000000001",--9587
"001111001100000010000000000000000001",--9588
"010110010001000001110000000000000111",--9589
"001111001010000001110000000000000010",--9590
"111110001100001001110011100000000000",--9591
"111110001110000001010011100000000001",--9592
"001111001100000010000000000000000010",--9593
"010110010001000001110000000000000010",--9594
"001011000000000001100000000100101111",--9595
"000101000000000000000010011001000001",--9596
"001111001010000001100000000000000001",--9597
"010010001101000000000000000000011001",--9598
"001101001000000001100000000000000100",--9599
"001101001000000001110000000000000110",--9600
"011010001101000000000000000000000010",--9601
"101001000000000010000000000000000001",--9602
"000101000000000000000010010110000101",--9603
"101000000001111000000100000000000000",--9604
"001111001100000001100000000000000001",--9605
"011100001111000010000000000000000001",--9606
"101110001101111000000011000000000010",--9607
"111110001100010001000011000000000000",--9608
"001111001010000001110000000000000001",--9609
"111110001110011000000011100000000000",--9610
"111110001100001001110011000000000000",--9611
"001111001010000001110000000000000010",--9612
"111110001100001001110011100000000000",--9613
"111110001110000001010011100000000001",--9614
"001111001100000010000000000000000010",--9615
"010110010001000001110000000000000111",--9616
"001111001010000001110000000000000000",--9617
"111110001100001001110011100000000000",--9618
"111110001110000000110011100000000001",--9619
"001111001100000010000000000000000000",--9620
"010110010001000001110000000000000010",--9621
"001011000000000001100000000100101111",--9622
"000101000000000000000010011001000001",--9623
"001111001010000001100000000000000010",--9624
"010010001101000000000000000111111010",--9625
"001101001000000001100000000000000100",--9626
"001101001000000001000000000000000110",--9627
"011010001101000000000000000000000010",--9628
"101001000000000001110000000000000001",--9629
"000101000000000000000010010110100000",--9630
"101000000001111000000011100000000000",--9631
"001111001100000001100000000000000010",--9632
"011100001001000001110000000000000001",--9633
"101110001101111000000011000000000010",--9634
"111110001100010001010010100000000000",--9635
"001111001010000001100000000000000010",--9636
"111110001100011000000011000000000000",--9637
"111110001010001001100010100000000000",--9638
"001111001010000001100000000000000000",--9639
"111110001010001001100011000000000000",--9640
"111110001100000000110001100000000001",--9641
"001111001100000001100000000000000000",--9642
"010110001101000000110000000111101000",--9643
"001111001010000000110000000000000001",--9644
"111110001010001000110001100000000000",--9645
"111110000110000001000001100000000001",--9646
"001111001100000001000000000000000001",--9647
"010110001001000000110000000111100011",--9648
"001011000000000001010000000100101111",--9649
"000101000000000000000010011001000001",--9650
"011111001011000000100000000000011010",--9651
"001101001000000001000000000000000100",--9652
"001101111100000001010000000000000000",--9653
"001111001010000001100000000000000000",--9654
"001111001000000001110000000000000000",--9655
"111110001100001001110011000000000000",--9656
"001111001010000001110000000000000001",--9657
"001111001000000010000000000000000001",--9658
"111110001110001010000011100000000000",--9659
"111110001100000001110011000000000000",--9660
"001111001010000001110000000000000010",--9661
"001111001000000010000000000000000010",--9662
"111110001110001010000011100000000000",--9663
"111110001100000001110011000000000000",--9664
"010110001101000000000000000111010010",--9665
"001111001000000001110000000000000000",--9666
"111110001110001000110001100000000000",--9667
"001111001000000001110000000000000001",--9668
"111110001110001001000010000000000000",--9669
"111110000110000001000001100000000000",--9670
"001111001000000001000000000000000010",--9671
"111110001000001001010010000000000000",--9672
"111110000110000001000001100000000010",--9673
"111110001100011000000010000000000000",--9674
"111110000110001001000001100000000000",--9675
"001011000000000000110000000100101111",--9676
"000101000000000000000010011001000001",--9677
"001101111100000001100000000000000000",--9678
"001111001100000001100000000000000000",--9679
"001111001100000001110000000000000001",--9680
"001111001100000010000000000000000010",--9681
"111110001100001001100100100000000000",--9682
"001101001000000001110000000000000100",--9683
"001111001110000010100000000000000000",--9684
"111110010010001010100100100000000000",--9685
"111110001110001001110101000000000000",--9686
"001111001110000010110000000000000001",--9687
"111110010100001010110101000000000000",--9688
"111110010010000010100100100000000000",--9689
"111110010000001010000101000000000000",--9690
"001111001110000010110000000000000010",--9691
"111110010100001010110101000000000000",--9692
"111110010010000010100100100000000000",--9693
"001101001000000010000000000000000011",--9694
"011100010001000000000000000000000011",--9695
"101110010011111000000011000000000000",--9696
"011110010011000000000000000000001111",--9697
"000101000000000000000010011110010100",--9698
"111110001110001010000101000000000000",--9699
"001101001000000010010000000000001001",--9700
"001111010010000010110000000000000000",--9701
"111110010100001010110101000000000000",--9702
"111110010010000010100100100000000000",--9703
"111110010000001001100100000000000000",--9704
"001111010010000010100000000000000001",--9705
"111110010000001010100100000000000000",--9706
"111110010010000010000100000000000000",--9707
"111110001100001001110011000000000000",--9708
"001111010010000001110000000000000010",--9709
"111110001100001001110011000000000000",--9710
"111110010000000001100011000000000000",--9711
"010010001101000000000000000110100011",--9712
"001111001100000001110000000000000000",--9713
"001111001100000010000000000000000001",--9714
"001111001100000010010000000000000010",--9715
"111110001110001000110101000000000000",--9716
"001111001110000010110000000000000000",--9717
"111110010100001010110101000000000000",--9718
"111110010000001001000101100000000000",--9719
"001111001110000011000000000000000001",--9720
"111110010110001011000101100000000000",--9721
"111110010100000010110101000000000000",--9722
"111110010010001001010101100000000000",--9723
"001111001110000011000000000000000010",--9724
"111110010110001011000101100000000000",--9725
"111110010100000010110101000000000000",--9726
"011100010001000000000000000000000010",--9727
"101110010101111000000011100000000000",--9728
"000101000000000000000010011000010111",--9729
"111110010010001001000101100000000000",--9730
"111110010000001001010110000000000000",--9731
"111110010110000011000101100000000000",--9732
"001101001000000010010000000000001001",--9733
"001111010010000011000000000000000000",--9734
"111110010110001011000101100000000000",--9735
"111110001110001001010110000000000000",--9736
"111110010010001000110100100000000000",--9737
"111110011000000010010100100000000000",--9738
"001111010010000011000000000000000001",--9739
"111110010010001011000100100000000000",--9740
"111110010110000010010100100000000000",--9741
"111110001110001001000011100000000000",--9742
"111110010000001000110100000000000000",--9743
"111110001110000010000011100000000000",--9744
"001111010010000010000000000000000010",--9745
"111110001110001010000011100000000000",--9746
"111110010010000001110011100000000000",--9747
"101111000001110010000011111100000000",--9748
"111110001110001010000011100000000000",--9749
"111110010100000001110011100000000000",--9750
"111110000110001000110100000000000000",--9751
"001111001110000010010000000000000000",--9752
"111110010000001010010100000000000000",--9753
"111110001000001001000100100000000000",--9754
"001111001110000010100000000000000001",--9755
"111110010010001010100100100000000000",--9756
"111110010000000010010100000000000000",--9757
"111110001010001001010100100000000000",--9758
"001111001110000010100000000000000010",--9759
"111110010010001010100100100000000000",--9760
"111110010000000010010100000000000000",--9761
"011100010001000000000000000000000011",--9762
"101110010001111000000001100000000000",--9763
"011111001011000000110000000000010000",--9764
"000101000000000000000010011000110100",--9765
"111110001000001001010100100000000000",--9766
"001101001000000001110000000000001001",--9767
"001111001110000010100000000000000000",--9768
"111110010010001010100100100000000000",--9769
"111110010000000010010100000000000000",--9770
"111110001010001000110010100000000000",--9771
"001111001110000010010000000000000001",--9772
"111110001010001010010010100000000000",--9773
"111110010000000001010010100000000000",--9774
"111110000110001001000001100000000000",--9775
"001111001110000001000000000000000010",--9776
"111110000110001001000001100000000000",--9777
"111110001010000000110001100000000000",--9778
"011111001011000000110000000000000001",--9779
"111110000110010000010001100000000000",--9780
"111110001110001001110010000000000000",--9781
"111110001100001000110001100000000000",--9782
"111110001000010000110001100000000000",--9783
"010110000111000000000000000101011011",--9784
"111110000110100000000001100000000000",--9785
"001101001000000001000000000000000110",--9786
"011100001001000000000000000000000001",--9787
"101110000111111000000001100000000010",--9788
"111110000110010001110001100000000000",--9789
"111110001100011000000010000000000000",--9790
"111110000110001001000001100000000000",--9791
"001011000000000000110000000100101111",--9792
"001111000000000000110000000100101111",--9793
"001111000000000001000000000100101101",--9794
"010110001001000000110000000101010000",--9795
"001101000100000001000000000000000001",--9796
"010011001001000000000000000101001110",--9797
"001101001000000001000000000100110001",--9798
"001101001000000001010000000000000000",--9799
"001001111100000000101111111111111100",--9800
"010011001011000000000000000100111001",--9801
"001101001010000001100000000101101101",--9802
"001111000000000000110000000100010101",--9803
"001101001100000001110000000000000101",--9804
"001111001110000001000000000000000000",--9805
"111110000110010001000001100000000000",--9806
"001111000000000001000000000100010110",--9807
"001111001110000001010000000000000001",--9808
"111110001000010001010010000000000000",--9809
"001111000000000001010000000100010111",--9810
"001111001110000001100000000000000010",--9811
"111110001010010001100010100000000000",--9812
"001101001100000001110000000000000001",--9813
"011111001111000000010000000001010101",--9814
"001101111100000001110000000000000000",--9815
"001111001110000001100000000000000000",--9816
"010010001101000000000000000000011010",--9817
"001101001100000010000000000000000100",--9818
"001101001100000010010000000000000110",--9819
"011010001101000000000000000000000010",--9820
"101001000000000010100000000000000001",--9821
"000101000000000000000010011001100000",--9822
"101000000001111000000101000000000000",--9823
"001111010000000001100000000000000000",--9824
"011100010011000010100000000000000001",--9825
"101110001101111000000011000000000010",--9826
"111110001100010000110011000000000000",--9827
"001111001110000001110000000000000000",--9828
"111110001110011000000011100000000000",--9829
"111110001100001001110011000000000000",--9830
"001111001110000001110000000000000001",--9831
"111110001100001001110011100000000000",--9832
"111110001110000001000011100000000001",--9833
"001111010000000010000000000000000001",--9834
"010110010001000001110000000000001000",--9835
"001111001110000001110000000000000010",--9836
"111110001100001001110011100000000000",--9837
"111110001110000001010011100000000001",--9838
"001111010000000010000000000000000010",--9839
"010110010001000001110000000000000011",--9840
"001011000000000001100000000100101111",--9841
"101001000000000001100000000000000001",--9842
"000101000000000000000010011101001001",--9843
"001111001110000001100000000000000001",--9844
"010010001101000000000000000000011010",--9845
"001101001100000010000000000000000100",--9846
"001101001100000010010000000000000110",--9847
"011010001101000000000000000000000010",--9848
"101001000000000010100000000000000001",--9849
"000101000000000000000010011001111100",--9850
"101000000001111000000101000000000000",--9851
"001111010000000001100000000000000001",--9852
"011100010011000010100000000000000001",--9853
"101110001101111000000011000000000010",--9854
"111110001100010001000011000000000000",--9855
"001111001110000001110000000000000001",--9856
"111110001110011000000011100000000000",--9857
"111110001100001001110011000000000000",--9858
"001111001110000001110000000000000010",--9859
"111110001100001001110011100000000000",--9860
"111110001110000001010011100000000001",--9861
"001111010000000010000000000000000010",--9862
"010110010001000001110000000000001000",--9863
"001111001110000001110000000000000000",--9864
"111110001100001001110011100000000000",--9865
"111110001110000000110011100000000001",--9866
"001111010000000010000000000000000000",--9867
"010110010001000001110000000000000011",--9868
"001011000000000001100000000100101111",--9869
"101001000000000001100000000000000010",--9870
"000101000000000000000010011101001001",--9871
"001111001110000001100000000000000010",--9872
"010010001101000000000000000010101011",--9873
"001101001100000010000000000000000100",--9874
"001101001100000001100000000000000110",--9875
"011010001101000000000000000000000010",--9876
"101001000000000010010000000000000001",--9877
"000101000000000000000010011010011000",--9878
"101000000001111000000100100000000000",--9879
"001111010000000001100000000000000010",--9880
"011100001101000010010000000000000001",--9881
"101110001101111000000011000000000010",--9882
"111110001100010001010010100000000000",--9883
"001111001110000001100000000000000010",--9884
"111110001100011000000011000000000000",--9885
"111110001010001001100010100000000000",--9886
"001111001110000001100000000000000000",--9887
"111110001010001001100011000000000000",--9888
"111110001100000000110001100000000001",--9889
"001111010000000001100000000000000000",--9890
"010110001101000000110000000010011001",--9891
"001111001110000000110000000000000001",--9892
"111110001010001000110001100000000000",--9893
"111110000110000001000001100000000001",--9894
"001111010000000001000000000000000001",--9895
"010110001001000000110000000010010100",--9896
"001011000000000001010000000100101111",--9897
"101001000000000001100000000000000011",--9898
"000101000000000000000010011101001001",--9899
"011111001111000000100000000000011011",--9900
"001101001100000001100000000000000100",--9901
"001101111100000001110000000000000000",--9902
"001111001110000001100000000000000000",--9903
"001111001100000001110000000000000000",--9904
"111110001100001001110011000000000000",--9905
"001111001110000001110000000000000001",--9906
"001111001100000010000000000000000001",--9907
"111110001110001010000011100000000000",--9908
"111110001100000001110011000000000000",--9909
"001111001110000001110000000000000010",--9910
"001111001100000010000000000000000010",--9911
"111110001110001010000011100000000000",--9912
"111110001100000001110011000000000000",--9913
"010110001101000000000000000010000010",--9914
"001111001100000001110000000000000000",--9915
"111110001110001000110001100000000000",--9916
"001111001100000001110000000000000001",--9917
"111110001110001001000010000000000000",--9918
"111110000110000001000001100000000000",--9919
"001111001100000001000000000000000010",--9920
"111110001000001001010010000000000000",--9921
"111110000110000001000001100000000010",--9922
"111110001100011000000010000000000000",--9923
"111110000110001001000001100000000000",--9924
"001011000000000000110000000100101111",--9925
"101001000000000001100000000000000001",--9926
"000101000000000000000010011101001001",--9927
"001101111100000010000000000000000000",--9928
"001111010000000001100000000000000000",--9929
"001111010000000001110000000000000001",--9930
"001111010000000010000000000000000010",--9931
"111110001100001001100100100000000000",--9932
"001101001100000010010000000000000100",--9933
"001111010010000010100000000000000000",--9934
"111110010010001010100100100000000000",--9935
"111110001110001001110101000000000000",--9936
"001111010010000010110000000000000001",--9937
"111110010100001010110101000000000000",--9938
"111110010010000010100100100000000000",--9939
"111110010000001010000101000000000000",--9940
"001111010010000010110000000000000010",--9941
"111110010100001010110101000000000000",--9942
"111110010010000010100100100000000000",--9943
"001101001100000010100000000000000011",--9944
"011100010101000000000000000000000011",--9945
"101110010011111000000011000000000000",--9946
"011110010011000000000000000000001111",--9947
"000101000000000000000010011100111101",--9948
"111110001110001010000101000000000000",--9949
"001101001100000010110000000000001001",--9950
"001111010110000010110000000000000000",--9951
"111110010100001010110101000000000000",--9952
"111110010010000010100100100000000000",--9953
"111110010000001001100100000000000000",--9954
"001111010110000010100000000000000001",--9955
"111110010000001010100100000000000000",--9956
"111110010010000010000100000000000000",--9957
"111110001100001001110011000000000000",--9958
"001111010110000001110000000000000010",--9959
"111110001100001001110011000000000000",--9960
"111110010000000001100011000000000000",--9961
"010010001101000000000000000001010010",--9962
"001111010000000001110000000000000000",--9963
"001111010000000010000000000000000001",--9964
"001111010000000010010000000000000010",--9965
"111110001110001000110101000000000000",--9966
"001111010010000010110000000000000000",--9967
"111110010100001010110101000000000000",--9968
"111110010000001001000101100000000000",--9969
"001111010010000011000000000000000001",--9970
"111110010110001011000101100000000000",--9971
"111110010100000010110101000000000000",--9972
"111110010010001001010101100000000000",--9973
"001111010010000011000000000000000010",--9974
"111110010110001011000101100000000000",--9975
"111110010100000010110101000000000000",--9976
"011100010101000000000000000000000010",--9977
"101110010101111000000011100000000000",--9978
"000101000000000000000010011100010001",--9979
"111110010010001001000101100000000000",--9980
"111110010000001001010110000000000000",--9981
"111110010110000011000101100000000000",--9982
"001101001100000010110000000000001001",--9983
"001111010110000011000000000000000000",--9984
"111110010110001011000101100000000000",--9985
"111110001110001001010110000000000000",--9986
"111110010010001000110100100000000000",--9987
"111110011000000010010100100000000000",--9988
"001111010110000011000000000000000001",--9989
"111110010010001011000100100000000000",--9990
"111110010110000010010100100000000000",--9991
"111110001110001001000011100000000000",--9992
"111110010000001000110100000000000000",--9993
"111110001110000010000011100000000000",--9994
"001111010110000010000000000000000010",--9995
"111110001110001010000011100000000000",--9996
"111110010010000001110011100000000000",--9997
"101111000001110010000011111100000000",--9998
"111110001110001010000011100000000000",--9999
"111110010100000001110011100000000000",--10000
"111110000110001000110100000000000000",--10001
"001111010010000010010000000000000000",--10002
"111110010000001010010100000000000000",--10003
"111110001000001001000100100000000000",--10004
"001111010010000010100000000000000001",--10005
"111110010010001010100100100000000000",--10006
"111110010000000010010100000000000000",--10007
"111110001010001001010100100000000000",--10008
"001111010010000010100000000000000010",--10009
"111110010010001010100100100000000000",--10010
"111110010000000010010100000000000000",--10011
"011100010101000000000000000000000011",--10012
"101110010001111000000001100000000000",--10013
"011111001111000000110000000000010000",--10014
"000101000000000000000010011100101110",--10015
"111110001000001001010100100000000000",--10016
"001101001100000010010000000000001001",--10017
"001111010010000010100000000000000000",--10018
"111110010010001010100100100000000000",--10019
"111110010000000010010100000000000000",--10020
"111110001010001000110010100000000000",--10021
"001111010010000010010000000000000001",--10022
"111110001010001010010010100000000000",--10023
"111110010000000001010010100000000000",--10024
"111110000110001001000001100000000000",--10025
"001111010010000001000000000000000010",--10026
"111110000110001001000001100000000000",--10027
"111110001010000000110001100000000000",--10028
"011111001111000000110000000000000001",--10029
"111110000110010000010001100000000000",--10030
"111110001110001001110010000000000000",--10031
"111110001100001000110001100000000000",--10032
"111110001000010000110001100000000000",--10033
"010110000111000000000000000000001010",--10034
"111110000110100000000001100000000000",--10035
"001101001100000001100000000000000110",--10036
"011100001101000000000000000000000001",--10037
"101110000111111000000001100000000010",--10038
"111110000110010001110001100000000000",--10039
"111110001100011000000010000000000000",--10040
"111110000110001001000001100000000000",--10041
"001011000000000000110000000100101111",--10042
"101001000000000001100000000000000001",--10043
"000101000000000000000010011101001001",--10044
"001101001010000001010000000101101101",--10045
"001101001010000001010000000000000110",--10046
"010000001011000000000000000001000011",--10047
"001101111100000000110000000000000000",--10048
"101000001001111000000001000000000000",--10049
"101001000000000000010000000000000001",--10050
"001001111100000111111111111111111011",--10051
"101001111100010111100000000000000110",--10052
"000111000000000000000001011101010010",--10053
"101001111100000111100000000000000110",--10054
"001101111100000111111111111111111011",--10055
"000101000000000000000010011110000011",--10056
"001111000000000000110000000100101111",--10057
"001001111100000001001111111111111011",--10058
"010110000111000000000000000000101111",--10059
"001111000000000001000000000100101101",--10060
"010110001001000000110000000000101101",--10061
"101111001001110001000011110000100011",--10062
"101111001001100001001101011100001010",--10063
"111110000110000001000001100000000000",--10064
"001101111100000001110000000000000000",--10065
"001111001110000001000000000000000000",--10066
"111110001000001000110010000000000000",--10067
"001111000000000001010000000100010101",--10068
"111110001000000001010010000000000000",--10069
"001111001110000001010000000000000001",--10070
"111110001010001000110010100000000000",--10071
"001111000000000001100000000100010110",--10072
"111110001010000001100010100000000000",--10073
"001111001110000001100000000000000010",--10074
"111110001100001000110011000000000000",--10075
"001111000000000001110000000100010111",--10076
"111110001100000001110011000000000000",--10077
"001001111100000001101111111111111010",--10078
"001001111100000001011111111111111001",--10079
"001011111100000001101111111111111000",--10080
"001011111100000001011111111111110111",--10081
"001011111100000001001111111111110110",--10082
"001011111100000000111111111111110101",--10083
"101000001001111000000001000000000000",--10084
"101000000001111000000000100000000000",--10085
"101110001001111000000001100000000000",--10086
"101110001011111000000010000000000000",--10087
"101110001101111000000010100000000000",--10088
"001001111100000111111111111111110100",--10089
"101001111100010111100000000000001101",--10090
"000111000000000000000000011110001000",--10091
"101001111100000111100000000000001101",--10092
"001101111100000111111111111111110100",--10093
"010000000011000000000000000000001100",--10094
"001111111100000000111111111111110101",--10095
"001011000000000000110000000100101101",--10096
"001111111100000000111111111111110110",--10097
"001011000000000000110000000100101010",--10098
"001111111100000000111111111111110111",--10099
"001011000000000000110000000100101011",--10100
"001111111100000000111111111111111000",--10101
"001011000000000000110000000100101100",--10102
"001101111100000000011111111111111001",--10103
"001001000000000000010000000100101001",--10104
"001101111100000000011111111111111010",--10105
"001001000000000000010000000100101110",--10106
"101001000000000000010000000000000001",--10107
"001101111100000000101111111111111011",--10108
"001101111100000000110000000000000000",--10109
"001001111100000111111111111111111010",--10110
"101001111100010111100000000000000111",--10111
"000111000000000000000001011101010010",--10112
"101001111100000111100000000000000111",--10113
"001101111100000111111111111111111010",--10114
"001101111100000000011111111111111100",--10115
"001101000010000000100000000000000010",--10116
"010011000101000000000000000000001110",--10117
"001101000100000000100000000100110001",--10118
"001101111100000000110000000000000000",--10119
"101000000001111000000000100000000000",--10120
"001001111100000111111111111111111011",--10121
"101001111100010111100000000000000110",--10122
"000111000000000000000001011101010010",--10123
"101001111100000111100000000000000110",--10124
"101001000000000000010000000000000011",--10125
"001101111100000000101111111111111100",--10126
"001101111100000000110000000000000000",--10127
"101001111100010111100000000000000110",--10128
"000111000000000000000001110100010111",--10129
"101001111100000111100000000000000110",--10130
"001101111100000111111111111111111011",--10131
"001101111100000000011111111111111101",--10132
"101001000010000000010000000000000001",--10133
"001101111100000000101111111111111111",--10134
"001101111100000000110000000000000000",--10135
"000101000000000000000010000001010110",--10136
"001100000100000000010010000000000000",--10137
"010011001000000000001111100000000000",--10138
"001101001000000001010000000101101101",--10139
"001101001010000001100000000000001010",--10140
"001111001100000000110000000000000000",--10141
"001111001100000001000000000000000001",--10142
"001111001100000001010000000000000010",--10143
"001101000110000001110000000000000001",--10144
"001100001110000001000100000000000000",--10145
"001101001010000010010000000000000001",--10146
"011111010011000000010000000000111011",--10147
"001101000110000001100000000000000000",--10148
"001111010000000001100000000000000000",--10149
"111110001100010000110011000000000000",--10150
"001111010000000001110000000000000001",--10151
"111110001100001001110011000000000000",--10152
"001111001100000001110000000000000001",--10153
"111110001100001001110011100000000000",--10154
"111110001110000001000011100000000001",--10155
"001101001010000001010000000000000100",--10156
"001111001010000010000000000000000001",--10157
"010110010001000001110000000000000111",--10158
"001111001100000001110000000000000010",--10159
"111110001100001001110011100000000000",--10160
"111110001110000001010011100000000001",--10161
"001111001010000010000000000000000010",--10162
"010110010001000001110000000000000010",--10163
"001111010000000001110000000000000001",--10164
"011110001111000000000000000000100110",--10165
"001111010000000001100000000000000010",--10166
"111110001100010001000011000000000000",--10167
"001111010000000001110000000000000011",--10168
"111110001100001001110011000000000000",--10169
"001111001100000001110000000000000000",--10170
"111110001100001001110011100000000000",--10171
"111110001110000000110011100000000001",--10172
"001111001010000010000000000000000000",--10173
"010110010001000001110000000000000111",--10174
"001111001100000001110000000000000010",--10175
"111110001100001001110011100000000000",--10176
"111110001110000001010011100000000001",--10177
"001111001010000010000000000000000010",--10178
"010110010001000001110000000000000010",--10179
"001111010000000001110000000000000011",--10180
"011110001111000000000000000000010011",--10181
"001111010000000001100000000000000100",--10182
"111110001100010001010010100000000000",--10183
"001111010000000001100000000000000101",--10184
"111110001010001001100010100000000000",--10185
"001111001100000001100000000000000000",--10186
"111110001010001001100011000000000000",--10187
"111110001100000000110001100000000001",--10188
"001111001010000001100000000000000000",--10189
"010110001101000000110000000000110110",--10190
"001111001100000000110000000000000001",--10191
"111110001010001000110001100000000000",--10192
"111110000110000001000001100000000001",--10193
"001111001010000001000000000000000001",--10194
"010110001001000000110000000000110001",--10195
"001111010000000000110000000000000101",--10196
"010010000111000000000000000000101111",--10197
"001011000000000001010000000100101111",--10198
"101001000000000001010000000000000011",--10199
"000101000000000000000010100101010011",--10200
"001011000000000001100000000100101111",--10201
"101001000000000001010000000000000010",--10202
"000101000000000000000010100101010011",--10203
"001011000000000001100000000100101111",--10204
"101001000000000001010000000000000001",--10205
"000101000000000000000010100101010011",--10206
"011111010011000000100000000000000111",--10207
"001111010000000000110000000000000000",--10208
"011010000111000000000000000000100011",--10209
"001111001100000001000000000000000011",--10210
"111110000110001001000001100000000000",--10211
"001011000000000000110000000100101111",--10212
"101001000000000001010000000000000001",--10213
"000101000000000000000010100101010011",--10214
"001111010000000001100000000000000000",--10215
"010010001101000000000000000000011100",--10216
"001111010000000001110000000000000001",--10217
"111110001110001000110001100000000000",--10218
"001111010000000001110000000000000010",--10219
"111110001110001001000010000000000000",--10220
"111110000110000001000001100000000000",--10221
"001111010000000001000000000000000011",--10222
"111110001000001001010010000000000000",--10223
"111110000110000001000001100000000000",--10224
"001111001100000001000000000000000011",--10225
"111110000110001000110010100000000000",--10226
"111110001100001001000010000000000000",--10227
"111110001010010001000010000000000000",--10228
"010110001001000000000000000000001111",--10229
"001101001010000001010000000000000110",--10230
"011100001011000000000000000000000110",--10231
"111110001000100000000010000000000000",--10232
"111110000110010001000001100000000000",--10233
"001111010000000001000000000000000100",--10234
"111110000110001001000001100000000000",--10235
"001011000000000000110000000100101111",--10236
"000101000000000000000010100000000011",--10237
"111110001000100000000010000000000000",--10238
"111110000110000001000001100000000000",--10239
"001111010000000001000000000000000100",--10240
"111110000110001001000001100000000000",--10241
"001011000000000000110000000100101111",--10242
"101001000000000001010000000000000001",--10243
"000101000000000000000010100101010011",--10244
"001101001000000001000000000101101101",--10245
"001101001000000001000000000000000110",--10246
"010000001000000000001111100000000000",--10247
"101001000010000000010000000000000001",--10248
"001100000100000000010010000000000000",--10249
"010011001000000000001111100000000000",--10250
"001101001000000001010000000101101101",--10251
"001101001010000001100000000000001010",--10252
"001111001100000000110000000000000000",--10253
"001111001100000001000000000000000001",--10254
"001111001100000001010000000000000010",--10255
"001100001110000001000011100000000000",--10256
"001101001010000010000000000000000001",--10257
"011111010001000000010000000000111011",--10258
"001101000110000001100000000000000000",--10259
"001111001110000001100000000000000000",--10260
"111110001100010000110011000000000000",--10261
"001111001110000001110000000000000001",--10262
"111110001100001001110011000000000000",--10263
"001111001100000001110000000000000001",--10264
"111110001100001001110011100000000000",--10265
"111110001110000001000011100000000001",--10266
"001101001010000001010000000000000100",--10267
"001111001010000010000000000000000001",--10268
"010110010001000001110000000000000111",--10269
"001111001100000001110000000000000010",--10270
"111110001100001001110011100000000000",--10271
"111110001110000001010011100000000001",--10272
"001111001010000010000000000000000010",--10273
"010110010001000001110000000000000010",--10274
"001111001110000001110000000000000001",--10275
"011110001111000000000000000000100110",--10276
"001111001110000001100000000000000010",--10277
"111110001100010001000011000000000000",--10278
"001111001110000001110000000000000011",--10279
"111110001100001001110011000000000000",--10280
"001111001100000001110000000000000000",--10281
"111110001100001001110011100000000000",--10282
"111110001110000000110011100000000001",--10283
"001111001010000010000000000000000000",--10284
"010110010001000001110000000000000111",--10285
"001111001100000001110000000000000010",--10286
"111110001100001001110011100000000000",--10287
"111110001110000001010011100000000001",--10288
"001111001010000010000000000000000010",--10289
"010110010001000001110000000000000010",--10290
"001111001110000001110000000000000011",--10291
"011110001111000000000000000000010011",--10292
"001111001110000001100000000000000100",--10293
"111110001100010001010010100000000000",--10294
"001111001110000001100000000000000101",--10295
"111110001010001001100010100000000000",--10296
"001111001100000001100000000000000000",--10297
"111110001010001001100011000000000000",--10298
"111110001100000000110001100000000001",--10299
"001111001010000001100000000000000000",--10300
"010110001101000000110000000000110110",--10301
"001111001100000000110000000000000001",--10302
"111110001010001000110001100000000000",--10303
"111110000110000001000001100000000001",--10304
"001111001010000001000000000000000001",--10305
"010110001001000000110000000000110001",--10306
"001111001110000000110000000000000101",--10307
"010010000111000000000000000000101111",--10308
"001011000000000001010000000100101111",--10309
"101001000000000001010000000000000011",--10310
"000101000000000000000010100001111001",--10311
"001011000000000001100000000100101111",--10312
"101001000000000001010000000000000010",--10313
"000101000000000000000010100001111001",--10314
"001011000000000001100000000100101111",--10315
"101001000000000001010000000000000001",--10316
"000101000000000000000010100001111001",--10317
"011111010001000000100000000000000111",--10318
"001111001110000000110000000000000000",--10319
"011010000111000000000000000000100011",--10320
"001111001100000001000000000000000011",--10321
"111110000110001001000001100000000000",--10322
"001011000000000000110000000100101111",--10323
"101001000000000001010000000000000001",--10324
"000101000000000000000010100001111001",--10325
"001111001110000001100000000000000000",--10326
"010010001101000000000000000000011100",--10327
"001111001110000001110000000000000001",--10328
"111110001110001000110001100000000000",--10329
"001111001110000001110000000000000010",--10330
"111110001110001001000010000000000000",--10331
"111110000110000001000001100000000000",--10332
"001111001110000001000000000000000011",--10333
"111110001000001001010010000000000000",--10334
"111110000110000001000001100000000000",--10335
"001111001100000001000000000000000011",--10336
"111110000110001000110010100000000000",--10337
"111110001100001001000010000000000000",--10338
"111110001010010001000010000000000000",--10339
"010110001001000000000000000000001111",--10340
"001101001010000001010000000000000110",--10341
"011100001011000000000000000000000110",--10342
"111110001000100000000010000000000000",--10343
"111110000110010001000001100000000000",--10344
"001111001110000001000000000000000100",--10345
"111110000110001001000001100000000000",--10346
"001011000000000000110000000100101111",--10347
"000101000000000000000010100001110010",--10348
"111110001000100000000010000000000000",--10349
"111110000110000001000001100000000000",--10350
"001111001110000001000000000000000100",--10351
"111110000110001001000001100000000000",--10352
"001011000000000000110000000100101111",--10353
"101001000000000001010000000000000001",--10354
"000101000000000000000010100001111001",--10355
"001101001000000001000000000101101101",--10356
"001101001000000001000000000000000110",--10357
"010000001000000000001111100000000000",--10358
"101001000010000000010000000000000001",--10359
"000101000000000000000010011110011001",--10360
"001111000000000000110000000100101111",--10361
"001001111100000000110000000000000000",--10362
"001001111100000000101111111111111111",--10363
"001001111100000000011111111111111110",--10364
"010110000111000000000000000011010000",--10365
"001111000000000001000000000100101101",--10366
"010110001001000000110000000011001110",--10367
"001101000110000001100000000000000000",--10368
"101111001001110001000011110000100011",--10369
"101111001001100001001101011100001010",--10370
"111110000110000001000001100000000000",--10371
"001111001100000001000000000000000000",--10372
"111110001000001000110010000000000000",--10373
"001111000000000001010000000100010010",--10374
"111110001000000001010010000000000000",--10375
"001111001100000001010000000000000001",--10376
"111110001010001000110010100000000000",--10377
"001111000000000001100000000100010011",--10378
"111110001010000001100010100000000000",--10379
"001111001100000001100000000000000010",--10380
"111110001100001000110011000000000000",--10381
"001111000000000001110000000100010100",--10382
"111110001100000001110011000000000000",--10383
"001101000100000001100000000000000000",--10384
"001001111100000001011111111111111101",--10385
"001001111100000001001111111111111100",--10386
"001011111100000001101111111111111011",--10387
"001011111100000001011111111111111010",--10388
"001011111100000001001111111111111001",--10389
"001011111100000000111111111111111000",--10390
"010011001101000000000000000010101010",--10391
"001101001100000001100000000101101101",--10392
"001101001100000001110000000000000101",--10393
"001111001110000001110000000000000000",--10394
"111110001000010001110011100000000000",--10395
"001111001110000010000000000000000001",--10396
"111110001010010010000100000000000000",--10397
"001111001110000010010000000000000010",--10398
"111110001100010010010100100000000000",--10399
"001101001100000001110000000000000001",--10400
"011111001111000000010000000000010000",--10401
"101110001111111000000011100000000001",--10402
"001101001100000001110000000000000100",--10403
"001111001110000010100000000000000000",--10404
"010110010101000001110000000000001001",--10405
"101110010001111000000011100000000001",--10406
"001111001110000010000000000000000001",--10407
"010110010001000001110000000000000110",--10408
"101110010011111000000011100000000001",--10409
"001111001110000010000000000000000010",--10410
"010110010001000001110000000000000011",--10411
"001101001100000001100000000000000110",--10412
"011100001101000000000000000010100000",--10413
"000101000000000000000010100011100111",--10414
"001101001100000001100000000000000110",--10415
"011100001101000000000000000000110110",--10416
"000101000000000000000010100101001110",--10417
"011111001111000000100000000000001111",--10418
"001101001100000001110000000000000100",--10419
"001111001110000010100000000000000000",--10420
"111110010100001001110011100000000000",--10421
"001111001110000010100000000000000001",--10422
"111110010100001010000100000000000000",--10423
"111110001110000010000011100000000000",--10424
"001111001110000010000000000000000010",--10425
"111110010000001010010100000000000000",--10426
"111110001110000010000011100000000000",--10427
"001101001100000001100000000000000110",--10428
"011010001111000000000000000000000010",--10429
"011111001101000000010000000000101000",--10430
"000101000000000000000010100101001110",--10431
"011100001101000000000000000000100110",--10432
"000101000000000000000010100101001110",--10433
"111110001110001001110101000000000000",--10434
"001101001100000010000000000000000100",--10435
"001111010000000010110000000000000000",--10436
"111110010100001010110101000000000000",--10437
"111110010000001010000101100000000000",--10438
"001111010000000011000000000000000001",--10439
"111110010110001011000101100000000000",--10440
"111110010100000010110101000000000000",--10441
"111110010010001010010101100000000000",--10442
"001111010000000011000000000000000010",--10443
"111110010110001011000101100000000000",--10444
"111110010100000010110101000000000000",--10445
"001101001100000010000000000000000011",--10446
"011100010001000000000000000000000011",--10447
"101110010101111000000011100000000000",--10448
"011111001111000000110000000000010000",--10449
"000101000000000000000010100011100001",--10450
"111110010000001010010101100000000000",--10451
"001101001100000010000000000000001001",--10452
"001111010000000011000000000000000000",--10453
"111110010110001011000101100000000000",--10454
"111110010100000010110101000000000000",--10455
"111110010010001001110100100000000000",--10456
"001111010000000010110000000000000001",--10457
"111110010010001010110100100000000000",--10458
"111110010100000010010100100000000000",--10459
"111110001110001010000011100000000000",--10460
"001111010000000010000000000000000010",--10461
"111110001110001010000011100000000000",--10462
"111110010010000001110011100000000000",--10463
"011111001111000000110000000000000001",--10464
"111110001110010000010011100000000000",--10465
"001101001100000001100000000000000110",--10466
"011010001111000000000000000000000010",--10467
"011111001101000000010000000000000010",--10468
"000101000000000000000010100101001110",--10469
"010000001101000000000000000001100111",--10470
"001101000100000001100000000000000001",--10471
"010011001101000000000000000001011001",--10472
"001101001100000001100000000101101101",--10473
"001101001100000001110000000000000101",--10474
"001111001110000001110000000000000000",--10475
"111110001000010001110011100000000000",--10476
"001111001110000010000000000000000001",--10477
"111110001010010010000100000000000000",--10478
"001111001110000010010000000000000010",--10479
"111110001100010010010100100000000000",--10480
"001101001100000001110000000000000001",--10481
"011111001111000000010000000000010000",--10482
"101110001111111000000011100000000001",--10483
"001101001100000001110000000000000100",--10484
"001111001110000010100000000000000000",--10485
"010110010101000001110000000000001001",--10486
"101110010001111000000011100000000001",--10487
"001111001110000010000000000000000001",--10488
"010110010001000001110000000000000110",--10489
"101110010011111000000011100000000001",--10490
"001111001110000010000000000000000010",--10491
"010110010001000001110000000000000011",--10492
"001101001100000001100000000000000110",--10493
"011100001101000000000000000001001111",--10494
"000101000000000000000010100100111000",--10495
"001101001100000001100000000000000110",--10496
"011100001101000000000000000000110110",--10497
"000101000000000000000010100101001110",--10498
"011111001111000000100000000000001111",--10499
"001101001100000001110000000000000100",--10500
"001111001110000010100000000000000000",--10501
"111110010100001001110011100000000000",--10502
"001111001110000010100000000000000001",--10503
"111110010100001010000100000000000000",--10504
"111110001110000010000011100000000000",--10505
"001111001110000010000000000000000010",--10506
"111110010000001010010100000000000000",--10507
"111110001110000010000011100000000000",--10508
"001101001100000001100000000000000110",--10509
"011010001111000000000000000000000010",--10510
"011111001101000000010000000000101000",--10511
"000101000000000000000010100101001110",--10512
"011100001101000000000000000000100110",--10513
"000101000000000000000010100101001110",--10514
"111110001110001001110101000000000000",--10515
"001101001100000010000000000000000100",--10516
"001111010000000010110000000000000000",--10517
"111110010100001010110101000000000000",--10518
"111110010000001010000101100000000000",--10519
"001111010000000011000000000000000001",--10520
"111110010110001011000101100000000000",--10521
"111110010100000010110101000000000000",--10522
"111110010010001010010101100000000000",--10523
"001111010000000011000000000000000010",--10524
"111110010110001011000101100000000000",--10525
"111110010100000010110101000000000000",--10526
"001101001100000010000000000000000011",--10527
"011100010001000000000000000000000011",--10528
"101110010101111000000011100000000000",--10529
"011111001111000000110000000000010000",--10530
"000101000000000000000010100100110010",--10531
"111110010000001010010101100000000000",--10532
"001101001100000010000000000000001001",--10533
"001111010000000011000000000000000000",--10534
"111110010110001011000101100000000000",--10535
"111110010100000010110101000000000000",--10536
"111110010010001001110100100000000000",--10537
"001111010000000010110000000000000001",--10538
"111110010010001010110100100000000000",--10539
"111110010100000010010100100000000000",--10540
"111110001110001010000011100000000000",--10541
"001111010000000010000000000000000010",--10542
"111110001110001010000011100000000000",--10543
"111110010010000001110011100000000000",--10544
"011111001111000000110000000000000001",--10545
"111110001110010000010011100000000000",--10546
"001101001100000001100000000000000110",--10547
"011010001111000000000000000000000010",--10548
"011111001101000000010000000000000010",--10549
"000101000000000000000010100101001110",--10550
"010000001101000000000000000000010110",--10551
"101001000000000000010000000000000010",--10552
"101110001001111000000001100000000000",--10553
"101110001011111000000010000000000000",--10554
"101110001101111000000010100000000000",--10555
"001001111100000111111111111111110111",--10556
"101001111100010111100000000000001010",--10557
"000111000000000000000000011110001000",--10558
"101001111100000111100000000000001010",--10559
"001101111100000111111111111111110111",--10560
"010000000011000000000000000000001100",--10561
"001111111100000000111111111111111000",--10562
"001011000000000000110000000100101101",--10563
"001111111100000000111111111111111001",--10564
"001011000000000000110000000100101010",--10565
"001111111100000000111111111111111010",--10566
"001011000000000000110000000100101011",--10567
"001111111100000000111111111111111011",--10568
"001011000000000000110000000100101100",--10569
"001101111100000000011111111111111100",--10570
"001001000000000000010000000100101001",--10571
"001101111100000000011111111111111101",--10572
"001001000000000000010000000100101110",--10573
"001101111100000000011111111111111110",--10574
"101001000010000000010000000000000001",--10575
"001101111100000000101111111111111111",--10576
"001101111100000000110000000000000000",--10577
"000101000000000000000010011110011001",--10578
"001111000000000000110000000100101111",--10579
"001001111100000000110000000000000000",--10580
"001001111100000001111111111111111111",--10581
"001001111100000000101111111111111110",--10582
"001001111100000000011111111111111101",--10583
"010110000111000000000000000100100001",--10584
"001111000000000001000000000100101101",--10585
"010110001001000000110000000100011111",--10586
"001101000110000001100000000000000000",--10587
"101111001001110001000011110000100011",--10588
"101111001001100001001101011100001010",--10589
"111110000110000001000001100000000000",--10590
"001111001100000001000000000000000000",--10591
"111110001000001000110010000000000000",--10592
"001111000000000001010000000100010010",--10593
"111110001000000001010010000000000000",--10594
"001111001100000001010000000000000001",--10595
"111110001010001000110010100000000000",--10596
"001111000000000001100000000100010011",--10597
"111110001010000001100010100000000000",--10598
"001111001100000001100000000000000010",--10599
"111110001100001000110011000000000000",--10600
"001111000000000001110000000100010100",--10601
"111110001100000001110011000000000000",--10602
"001101000100000001100000000000000000",--10603
"001001111100000001011111111111111100",--10604
"001001111100000001001111111111111011",--10605
"001011111100000001101111111111111010",--10606
"001011111100000001011111111111111001",--10607
"001011111100000001001111111111111000",--10608
"001011111100000000111111111111110111",--10609
"010011001101000000000000000011111011",--10610
"001101001100000001100000000101101101",--10611
"001101001100000010000000000000000101",--10612
"001111010000000001110000000000000000",--10613
"111110001000010001110011100000000000",--10614
"001111010000000010000000000000000001",--10615
"111110001010010010000100000000000000",--10616
"001111010000000010010000000000000010",--10617
"111110001100010010010100100000000000",--10618
"001101001100000010000000000000000001",--10619
"011111010001000000010000000000010000",--10620
"101110001111111000000011100000000001",--10621
"001101001100000010000000000000000100",--10622
"001111010000000010100000000000000000",--10623
"010110010101000001110000000000001001",--10624
"101110010001111000000011100000000001",--10625
"001111010000000010000000000000000001",--10626
"010110010001000001110000000000000110",--10627
"101110010011111000000011100000000001",--10628
"001111010000000010000000000000000010",--10629
"010110010001000001110000000000000011",--10630
"001101001100000001100000000000000110",--10631
"011100001101000000000000000011110001",--10632
"000101000000000000000010100111000010",--10633
"001101001100000001100000000000000110",--10634
"011100001101000000000000000000110110",--10635
"000101000000000000000010101001111010",--10636
"011111010001000000100000000000001111",--10637
"001101001100000010000000000000000100",--10638
"001111010000000010100000000000000000",--10639
"111110010100001001110011100000000000",--10640
"001111010000000010100000000000000001",--10641
"111110010100001010000100000000000000",--10642
"111110001110000010000011100000000000",--10643
"001111010000000010000000000000000010",--10644
"111110010000001010010100000000000000",--10645
"111110001110000010000011100000000000",--10646
"001101001100000001100000000000000110",--10647
"011010001111000000000000000000000010",--10648
"011111001101000000010000000000101000",--10649
"000101000000000000000010101001111010",--10650
"011100001101000000000000000000100110",--10651
"000101000000000000000010101001111010",--10652
"111110001110001001110101000000000000",--10653
"001101001100000010010000000000000100",--10654
"001111010010000010110000000000000000",--10655
"111110010100001010110101000000000000",--10656
"111110010000001010000101100000000000",--10657
"001111010010000011000000000000000001",--10658
"111110010110001011000101100000000000",--10659
"111110010100000010110101000000000000",--10660
"111110010010001010010101100000000000",--10661
"001111010010000011000000000000000010",--10662
"111110010110001011000101100000000000",--10663
"111110010100000010110101000000000000",--10664
"001101001100000010010000000000000011",--10665
"011100010011000000000000000000000011",--10666
"101110010101111000000011100000000000",--10667
"011111010001000000110000000000010000",--10668
"000101000000000000000010100110111100",--10669
"111110010000001010010101100000000000",--10670
"001101001100000010010000000000001001",--10671
"001111010010000011000000000000000000",--10672
"111110010110001011000101100000000000",--10673
"111110010100000010110101000000000000",--10674
"111110010010001001110100100000000000",--10675
"001111010010000010110000000000000001",--10676
"111110010010001010110100100000000000",--10677
"111110010100000010010100100000000000",--10678
"111110001110001010000011100000000000",--10679
"001111010010000010000000000000000010",--10680
"111110001110001010000011100000000000",--10681
"111110010010000001110011100000000000",--10682
"011111010001000000110000000000000001",--10683
"111110001110010000010011100000000000",--10684
"001101001100000001100000000000000110",--10685
"011010001111000000000000000000000010",--10686
"011111001101000000010000000000000010",--10687
"000101000000000000000010101001111010",--10688
"010000001101000000000000000010111000",--10689
"001101000100000001100000000000000001",--10690
"010011001101000000000000000010101010",--10691
"001101001100000001100000000101101101",--10692
"001101001100000010000000000000000101",--10693
"001111010000000001110000000000000000",--10694
"111110001000010001110011100000000000",--10695
"001111010000000010000000000000000001",--10696
"111110001010010010000100000000000000",--10697
"001111010000000010010000000000000010",--10698
"111110001100010010010100100000000000",--10699
"001101001100000010000000000000000001",--10700
"011111010001000000010000000000010000",--10701
"101110001111111000000011100000000001",--10702
"001101001100000010000000000000000100",--10703
"001111010000000010100000000000000000",--10704
"010110010101000001110000000000001001",--10705
"101110010001111000000011100000000001",--10706
"001111010000000010000000000000000001",--10707
"010110010001000001110000000000000110",--10708
"101110010011111000000011100000000001",--10709
"001111010000000010000000000000000010",--10710
"010110010001000001110000000000000011",--10711
"001101001100000001100000000000000110",--10712
"011100001101000000000000000010100000",--10713
"000101000000000000000010101000010011",--10714
"001101001100000001100000000000000110",--10715
"011100001101000000000000000000110110",--10716
"000101000000000000000010101001111010",--10717
"011111010001000000100000000000001111",--10718
"001101001100000010000000000000000100",--10719
"001111010000000010100000000000000000",--10720
"111110010100001001110011100000000000",--10721
"001111010000000010100000000000000001",--10722
"111110010100001010000100000000000000",--10723
"111110001110000010000011100000000000",--10724
"001111010000000010000000000000000010",--10725
"111110010000001010010100000000000000",--10726
"111110001110000010000011100000000000",--10727
"001101001100000001100000000000000110",--10728
"011010001111000000000000000000000010",--10729
"011111001101000000010000000000101000",--10730
"000101000000000000000010101001111010",--10731
"011100001101000000000000000000100110",--10732
"000101000000000000000010101001111010",--10733
"111110001110001001110101000000000000",--10734
"001101001100000010010000000000000100",--10735
"001111010010000010110000000000000000",--10736
"111110010100001010110101000000000000",--10737
"111110010000001010000101100000000000",--10738
"001111010010000011000000000000000001",--10739
"111110010110001011000101100000000000",--10740
"111110010100000010110101000000000000",--10741
"111110010010001010010101100000000000",--10742
"001111010010000011000000000000000010",--10743
"111110010110001011000101100000000000",--10744
"111110010100000010110101000000000000",--10745
"001101001100000010010000000000000011",--10746
"011100010011000000000000000000000011",--10747
"101110010101111000000011100000000000",--10748
"011111010001000000110000000000010000",--10749
"000101000000000000000010101000001101",--10750
"111110010000001010010101100000000000",--10751
"001101001100000010010000000000001001",--10752
"001111010010000011000000000000000000",--10753
"111110010110001011000101100000000000",--10754
"111110010100000010110101000000000000",--10755
"111110010010001001110100100000000000",--10756
"001111010010000010110000000000000001",--10757
"111110010010001010110100100000000000",--10758
"111110010100000010010100100000000000",--10759
"111110001110001010000011100000000000",--10760
"001111010010000010000000000000000010",--10761
"111110001110001010000011100000000000",--10762
"111110010010000001110011100000000000",--10763
"011111010001000000110000000000000001",--10764
"111110001110010000010011100000000000",--10765
"001101001100000001100000000000000110",--10766
"011010001111000000000000000000000010",--10767
"011111001101000000010000000000000010",--10768
"000101000000000000000010101001111010",--10769
"010000001101000000000000000001100111",--10770
"001101000100000001100000000000000010",--10771
"010011001101000000000000000001011001",--10772
"001101001100000001100000000101101101",--10773
"001101001100000010000000000000000101",--10774
"001111010000000001110000000000000000",--10775
"111110001000010001110011100000000000",--10776
"001111010000000010000000000000000001",--10777
"111110001010010010000100000000000000",--10778
"001111010000000010010000000000000010",--10779
"111110001100010010010100100000000000",--10780
"001101001100000010000000000000000001",--10781
"011111010001000000010000000000010000",--10782
"101110001111111000000011100000000001",--10783
"001101001100000010000000000000000100",--10784
"001111010000000010100000000000000000",--10785
"010110010101000001110000000000001001",--10786
"101110010001111000000011100000000001",--10787
"001111010000000010000000000000000001",--10788
"010110010001000001110000000000000110",--10789
"101110010011111000000011100000000001",--10790
"001111010000000010000000000000000010",--10791
"010110010001000001110000000000000011",--10792
"001101001100000001100000000000000110",--10793
"011100001101000000000000000001001111",--10794
"000101000000000000000010101001100100",--10795
"001101001100000001100000000000000110",--10796
"011100001101000000000000000000110110",--10797
"000101000000000000000010101001111010",--10798
"011111010001000000100000000000001111",--10799
"001101001100000010000000000000000100",--10800
"001111010000000010100000000000000000",--10801
"111110010100001001110011100000000000",--10802
"001111010000000010100000000000000001",--10803
"111110010100001010000100000000000000",--10804
"111110001110000010000011100000000000",--10805
"001111010000000010000000000000000010",--10806
"111110010000001010010100000000000000",--10807
"111110001110000010000011100000000000",--10808
"001101001100000001100000000000000110",--10809
"011010001111000000000000000000000010",--10810
"011111001101000000010000000000101000",--10811
"000101000000000000000010101001111010",--10812
"011100001101000000000000000000100110",--10813
"000101000000000000000010101001111010",--10814
"111110001110001001110101000000000000",--10815
"001101001100000010010000000000000100",--10816
"001111010010000010110000000000000000",--10817
"111110010100001010110101000000000000",--10818
"111110010000001010000101100000000000",--10819
"001111010010000011000000000000000001",--10820
"111110010110001011000101100000000000",--10821
"111110010100000010110101000000000000",--10822
"111110010010001010010101100000000000",--10823
"001111010010000011000000000000000010",--10824
"111110010110001011000101100000000000",--10825
"111110010100000010110101000000000000",--10826
"001101001100000010010000000000000011",--10827
"011100010011000000000000000000000011",--10828
"101110010101111000000011100000000000",--10829
"011111010001000000110000000000010000",--10830
"000101000000000000000010101001011110",--10831
"111110010000001010010101100000000000",--10832
"001101001100000010010000000000001001",--10833
"001111010010000011000000000000000000",--10834
"111110010110001011000101100000000000",--10835
"111110010100000010110101000000000000",--10836
"111110010010001001110100100000000000",--10837
"001111010010000010110000000000000001",--10838
"111110010010001010110100100000000000",--10839
"111110010100000010010100100000000000",--10840
"111110001110001010000011100000000000",--10841
"001111010010000010000000000000000010",--10842
"111110001110001010000011100000000000",--10843
"111110010010000001110011100000000000",--10844
"011111010001000000110000000000000001",--10845
"111110001110010000010011100000000000",--10846
"001101001100000001100000000000000110",--10847
"011010001111000000000000000000000010",--10848
"011111001101000000010000000000000010",--10849
"000101000000000000000010101001111010",--10850
"010000001101000000000000000000010110",--10851
"101001000000000000010000000000000011",--10852
"101110001001111000000001100000000000",--10853
"101110001011111000000010000000000000",--10854
"101110001101111000000010100000000000",--10855
"001001111100000111111111111111110110",--10856
"101001111100010111100000000000001011",--10857
"000111000000000000000000011110001000",--10858
"101001111100000111100000000000001011",--10859
"001101111100000111111111111111110110",--10860
"010000000011000000000000000000001100",--10861
"001111111100000000111111111111110111",--10862
"001011000000000000110000000100101101",--10863
"001111111100000000111111111111111000",--10864
"001011000000000000110000000100101010",--10865
"001111111100000000111111111111111001",--10866
"001011000000000000110000000100101011",--10867
"001111111100000000111111111111111010",--10868
"001011000000000000110000000100101100",--10869
"001101111100000000011111111111111011",--10870
"001001000000000000010000000100101001",--10871
"001101111100000000011111111111111100",--10872
"001001000000000000010000000100101110",--10873
"001101111100000000011111111111111101",--10874
"101001000010000000010000000000000001",--10875
"001101111100000000111111111111111110",--10876
"001100000110000000010001000000000000",--10877
"010011000100000000001111100000000000",--10878
"001101000100000001000000000101101101",--10879
"001101001000000001010000000000001010",--10880
"001111001010000000110000000000000000",--10881
"001111001010000001000000000000000001",--10882
"001111001010000001010000000000000010",--10883
"001101111100000001111111111111111111",--10884
"001100001110000000100011000000000000",--10885
"001101001000000001110000000000000001",--10886
"011111001111000000010000000000111100",--10887
"001101111100000001010000000000000000",--10888
"001101001010000001110000000000000000",--10889
"001111001100000001100000000000000000",--10890
"111110001100010000110011000000000000",--10891
"001111001100000001110000000000000001",--10892
"111110001100001001110011000000000000",--10893
"001111001110000001110000000000000001",--10894
"111110001100001001110011100000000000",--10895
"111110001110000001000011100000000001",--10896
"001101001000000001000000000000000100",--10897
"001111001000000010000000000000000001",--10898
"010110010001000001110000000000000111",--10899
"001111001110000001110000000000000010",--10900
"111110001100001001110011100000000000",--10901
"111110001110000001010011100000000001",--10902
"001111001000000010000000000000000010",--10903
"010110010001000001110000000000000010",--10904
"001111001100000001110000000000000001",--10905
"011110001111000000000000000000100110",--10906
"001111001100000001100000000000000010",--10907
"111110001100010001000011000000000000",--10908
"001111001100000001110000000000000011",--10909
"111110001100001001110011000000000000",--10910
"001111001110000001110000000000000000",--10911
"111110001100001001110011100000000000",--10912
"111110001110000000110011100000000001",--10913
"001111001000000010000000000000000000",--10914
"010110010001000001110000000000000111",--10915
"001111001110000001110000000000000010",--10916
"111110001100001001110011100000000000",--10917
"111110001110000001010011100000000001",--10918
"001111001000000010000000000000000010",--10919
"010110010001000001110000000000000010",--10920
"001111001100000001110000000000000011",--10921
"011110001111000000000000000000010011",--10922
"001111001100000001100000000000000100",--10923
"111110001100010001010010100000000000",--10924
"001111001100000001100000000000000101",--10925
"111110001010001001100010100000000000",--10926
"001111001110000001100000000000000000",--10927
"111110001010001001100011000000000000",--10928
"111110001100000000110001100000000001",--10929
"001111001000000001100000000000000000",--10930
"010110001101000000110000000000110110",--10931
"001111001110000000110000000000000001",--10932
"111110001010001000110001100000000000",--10933
"111110000110000001000001100000000001",--10934
"001111001000000001000000000000000001",--10935
"010110001001000000110000000000110001",--10936
"001111001100000000110000000000000101",--10937
"010010000111000000000000000000101111",--10938
"001011000000000001010000000100101111",--10939
"101001000000000001000000000000000011",--10940
"000101000000000000000010101011110011",--10941
"001011000000000001100000000100101111",--10942
"101001000000000001000000000000000010",--10943
"000101000000000000000010101011110011",--10944
"001011000000000001100000000100101111",--10945
"101001000000000001000000000000000001",--10946
"000101000000000000000010101011110011",--10947
"011111001111000000100000000000000111",--10948
"001111001100000000110000000000000000",--10949
"011010000111000000000000000000100011",--10950
"001111001010000001000000000000000011",--10951
"111110000110001001000001100000000000",--10952
"001011000000000000110000000100101111",--10953
"101001000000000001000000000000000001",--10954
"000101000000000000000010101011110011",--10955
"001111001100000001100000000000000000",--10956
"010010001101000000000000000000011100",--10957
"001111001100000001110000000000000001",--10958
"111110001110001000110001100000000000",--10959
"001111001100000001110000000000000010",--10960
"111110001110001001000010000000000000",--10961
"111110000110000001000001100000000000",--10962
"001111001100000001000000000000000011",--10963
"111110001000001001010010000000000000",--10964
"111110000110000001000001100000000000",--10965
"001111001010000001000000000000000011",--10966
"111110000110001000110010100000000000",--10967
"111110001100001001000010000000000000",--10968
"111110001010010001000010000000000000",--10969
"010110001001000000000000000000001111",--10970
"001101001000000001000000000000000110",--10971
"011100001001000000000000000000000110",--10972
"111110001000100000000010000000000000",--10973
"111110000110010001000001100000000000",--10974
"001111001100000001000000000000000100",--10975
"111110000110001001000001100000000000",--10976
"001011000000000000110000000100101111",--10977
"000101000000000000000010101011101000",--10978
"111110001000100000000010000000000000",--10979
"111110000110000001000001100000000000",--10980
"001111001100000001000000000000000100",--10981
"111110000110001001000001100000000000",--10982
"001011000000000000110000000100101111",--10983
"101001000000000001000000000000000001",--10984
"000101000000000000000010101011110011",--10985
"001101000100000000100000000101101101",--10986
"001101000100000000100000000000000110",--10987
"010000000100000000001111100000000000",--10988
"101001000010000000010000000000000001",--10989
"001101111100000000100000000000000000",--10990
"101000000111111000001101100000000000",--10991
"101000000101111000000001100000000000",--10992
"101000110111111000000001000000000000",--10993
"000101000000000000000010011110011001",--10994
"001111000000000000110000000100101111",--10995
"001001111100000000011111111111111100",--10996
"010110000111000000000000000011010010",--10997
"001111000000000001000000000100101101",--10998
"010110001001000000110000000011010000",--10999
"001101111100000001010000000000000000",--11000
"001101001010000001100000000000000000",--11001
"101111001001110001000011110000100011",--11002
"101111001001100001001101011100001010",--11003
"111110000110000001000001100000000000",--11004
"001111001100000001000000000000000000",--11005
"111110001000001000110010000000000000",--11006
"001111000000000001010000000100010010",--11007
"111110001000000001010010000000000000",--11008
"001111001100000001010000000000000001",--11009
"111110001010001000110010100000000000",--11010
"001111000000000001100000000100010011",--11011
"111110001010000001100010100000000000",--11012
"001111001100000001100000000000000010",--11013
"111110001100001000110011000000000000",--11014
"001111000000000001110000000100010100",--11015
"111110001100000001110011000000000000",--11016
"001101000110000001100000000000000000",--11017
"001001111100000001001111111111111011",--11018
"001001111100000000101111111111111010",--11019
"001011111100000001101111111111111001",--11020
"001011111100000001011111111111111000",--11021
"001011111100000001001111111111110111",--11022
"001011111100000000111111111111110110",--11023
"010011001101000000000000000010101011",--11024
"001101001100000001100000000101101101",--11025
"001101001100000001110000000000000101",--11026
"001111001110000001110000000000000000",--11027
"111110001000010001110011100000000000",--11028
"001111001110000010000000000000000001",--11029
"111110001010010010000100000000000000",--11030
"001111001110000010010000000000000010",--11031
"111110001100010010010100100000000000",--11032
"001101001100000001110000000000000001",--11033
"011111001111000000010000000000010000",--11034
"101110001111111000000011100000000001",--11035
"001101001100000001110000000000000100",--11036
"001111001110000010100000000000000000",--11037
"010110010101000001110000000000001001",--11038
"101110010001111000000011100000000001",--11039
"001111001110000010000000000000000001",--11040
"010110010001000001110000000000000110",--11041
"101110010011111000000011100000000001",--11042
"001111001110000010000000000000000010",--11043
"010110010001000001110000000000000011",--11044
"001101001100000001100000000000000110",--11045
"011100001101000000000000000010100001",--11046
"000101000000000000000010101101100000",--11047
"001101001100000001100000000000000110",--11048
"011100001101000000000000000000110110",--11049
"000101000000000000000010101111001000",--11050
"011111001111000000100000000000001111",--11051
"001101001100000001110000000000000100",--11052
"001111001110000010100000000000000000",--11053
"111110010100001001110011100000000000",--11054
"001111001110000010100000000000000001",--11055
"111110010100001010000100000000000000",--11056
"111110001110000010000011100000000000",--11057
"001111001110000010000000000000000010",--11058
"111110010000001010010100000000000000",--11059
"111110001110000010000011100000000000",--11060
"001101001100000001100000000000000110",--11061
"011010001111000000000000000000000010",--11062
"011111001101000000010000000000101000",--11063
"000101000000000000000010101111001000",--11064
"011100001101000000000000000000100110",--11065
"000101000000000000000010101111001000",--11066
"111110001110001001110101000000000000",--11067
"001101001100000010000000000000000100",--11068
"001111010000000010110000000000000000",--11069
"111110010100001010110101000000000000",--11070
"111110010000001010000101100000000000",--11071
"001111010000000011000000000000000001",--11072
"111110010110001011000101100000000000",--11073
"111110010100000010110101000000000000",--11074
"111110010010001010010101100000000000",--11075
"001111010000000011000000000000000010",--11076
"111110010110001011000101100000000000",--11077
"111110010100000010110101000000000000",--11078
"001101001100000010000000000000000011",--11079
"011100010001000000000000000000000011",--11080
"101110010101111000000011100000000000",--11081
"011111001111000000110000000000010000",--11082
"000101000000000000000010101101011010",--11083
"111110010000001010010101100000000000",--11084
"001101001100000010000000000000001001",--11085
"001111010000000011000000000000000000",--11086
"111110010110001011000101100000000000",--11087
"111110010100000010110101000000000000",--11088
"111110010010001001110100100000000000",--11089
"001111010000000010110000000000000001",--11090
"111110010010001010110100100000000000",--11091
"111110010100000010010100100000000000",--11092
"111110001110001010000011100000000000",--11093
"001111010000000010000000000000000010",--11094
"111110001110001010000011100000000000",--11095
"111110010010000001110011100000000000",--11096
"011111001111000000110000000000000001",--11097
"111110001110010000010011100000000000",--11098
"001101001100000001100000000000000110",--11099
"011010001111000000000000000000000010",--11100
"011111001101000000010000000000000010",--11101
"000101000000000000000010101111001000",--11102
"010000001101000000000000000001101000",--11103
"001101000110000001100000000000000001",--11104
"010011001101000000000000000001011010",--11105
"001101001100000001100000000101101101",--11106
"001101001100000001110000000000000101",--11107
"001111001110000001110000000000000000",--11108
"111110001000010001110011100000000000",--11109
"001111001110000010000000000000000001",--11110
"111110001010010010000100000000000000",--11111
"001111001110000010010000000000000010",--11112
"111110001100010010010100100000000000",--11113
"001101001100000001110000000000000001",--11114
"011111001111000000010000000000010000",--11115
"101110001111111000000011100000000001",--11116
"001101001100000001110000000000000100",--11117
"001111001110000010100000000000000000",--11118
"010110010101000001110000000000001001",--11119
"101110010001111000000011100000000001",--11120
"001111001110000010000000000000000001",--11121
"010110010001000001110000000000000110",--11122
"101110010011111000000011100000000001",--11123
"001111001110000010000000000000000010",--11124
"010110010001000001110000000000000011",--11125
"001101001100000001100000000000000110",--11126
"011100001101000000000000000001010000",--11127
"000101000000000000000010101110110001",--11128
"001101001100000001100000000000000110",--11129
"011100001101000000000000000000110110",--11130
"000101000000000000000010101111001000",--11131
"011111001111000000100000000000001111",--11132
"001101001100000001110000000000000100",--11133
"001111001110000010100000000000000000",--11134
"111110010100001001110011100000000000",--11135
"001111001110000010100000000000000001",--11136
"111110010100001010000100000000000000",--11137
"111110001110000010000011100000000000",--11138
"001111001110000010000000000000000010",--11139
"111110010000001010010100000000000000",--11140
"111110001110000010000011100000000000",--11141
"001101001100000001100000000000000110",--11142
"011010001111000000000000000000000010",--11143
"011111001101000000010000000000101000",--11144
"000101000000000000000010101111001000",--11145
"011100001101000000000000000000100110",--11146
"000101000000000000000010101111001000",--11147
"111110001110001001110101000000000000",--11148
"001101001100000010000000000000000100",--11149
"001111010000000010110000000000000000",--11150
"111110010100001010110101000000000000",--11151
"111110010000001010000101100000000000",--11152
"001111010000000011000000000000000001",--11153
"111110010110001011000101100000000000",--11154
"111110010100000010110101000000000000",--11155
"111110010010001010010101100000000000",--11156
"001111010000000011000000000000000010",--11157
"111110010110001011000101100000000000",--11158
"111110010100000010110101000000000000",--11159
"001101001100000010000000000000000011",--11160
"011100010001000000000000000000000011",--11161
"101110010101111000000011100000000000",--11162
"011111001111000000110000000000010000",--11163
"000101000000000000000010101110101011",--11164
"111110010000001010010101100000000000",--11165
"001101001100000010000000000000001001",--11166
"001111010000000011000000000000000000",--11167
"111110010110001011000101100000000000",--11168
"111110010100000010110101000000000000",--11169
"111110010010001001110100100000000000",--11170
"001111010000000010110000000000000001",--11171
"111110010010001010110100100000000000",--11172
"111110010100000010010100100000000000",--11173
"111110001110001010000011100000000000",--11174
"001111010000000010000000000000000010",--11175
"111110001110001010000011100000000000",--11176
"111110010010000001110011100000000000",--11177
"011111001111000000110000000000000001",--11178
"111110001110010000010011100000000000",--11179
"001101001100000001100000000000000110",--11180
"011010001111000000000000000000000010",--11181
"011111001101000000010000000000000010",--11182
"000101000000000000000010101111001000",--11183
"010000001101000000000000000000010111",--11184
"101000000111111000000001000000000000",--11185
"101001000000000000010000000000000010",--11186
"101110001001111000000001100000000000",--11187
"101110001011111000000010000000000000",--11188
"101110001101111000000010100000000000",--11189
"001001111100000111111111111111110101",--11190
"101001111100010111100000000000001100",--11191
"000111000000000000000000011110001000",--11192
"101001111100000111100000000000001100",--11193
"001101111100000111111111111111110101",--11194
"010000000011000000000000000000001100",--11195
"001111111100000000111111111111110110",--11196
"001011000000000000110000000100101101",--11197
"001111111100000000111111111111110111",--11198
"001011000000000000110000000100101010",--11199
"001111111100000000111111111111111000",--11200
"001011000000000000110000000100101011",--11201
"001111111100000000111111111111111001",--11202
"001011000000000000110000000100101100",--11203
"001101111100000000011111111111111010",--11204
"001001000000000000010000000100101001",--11205
"001101111100000000011111111111111011",--11206
"001001000000000000010000000100101110",--11207
"001101111100000000011111111111111100",--11208
"101001000010000000010000000000000001",--11209
"001101111100000000101111111111111110",--11210
"001101111100000000110000000000000000",--11211
"000101000000000000000010011110011001",--11212
"001100000100000000010010000000000000",--11213
"010011001000000000001111100000000000",--11214
"001101001000000001000000000100110001",--11215
"001101001000000001010000000000000000",--11216
"001001111100000000110000000000000000",--11217
"001001111100000000101111111111111111",--11218
"001001111100000000011111111111111110",--11219
"010011001011000000000000000101010001",--11220
"001101001010000001100000000101101101",--11221
"001101001100000001110000000000001010",--11222
"001111001110000000110000000000000000",--11223
"001111001110000001000000000000000001",--11224
"001111001110000001010000000000000010",--11225
"001101000110000010000000000000000001",--11226
"001100010000000001010100000000000000",--11227
"001101001100000010010000000000000001",--11228
"011111010011000000010000000000111011",--11229
"001101000110000001110000000000000000",--11230
"001111010000000001100000000000000000",--11231
"111110001100010000110011000000000000",--11232
"001111010000000001110000000000000001",--11233
"111110001100001001110011000000000000",--11234
"001111001110000001110000000000000001",--11235
"111110001100001001110011100000000000",--11236
"111110001110000001000011100000000001",--11237
"001101001100000001100000000000000100",--11238
"001111001100000010000000000000000001",--11239
"010110010001000001110000000000000111",--11240
"001111001110000001110000000000000010",--11241
"111110001100001001110011100000000000",--11242
"111110001110000001010011100000000001",--11243
"001111001100000010000000000000000010",--11244
"010110010001000001110000000000000010",--11245
"001111010000000001110000000000000001",--11246
"011110001111000000000000000000100110",--11247
"001111010000000001100000000000000010",--11248
"111110001100010001000011000000000000",--11249
"001111010000000001110000000000000011",--11250
"111110001100001001110011000000000000",--11251
"001111001110000001110000000000000000",--11252
"111110001100001001110011100000000000",--11253
"111110001110000000110011100000000001",--11254
"001111001100000010000000000000000000",--11255
"010110010001000001110000000000000111",--11256
"001111001110000001110000000000000010",--11257
"111110001100001001110011100000000000",--11258
"111110001110000001010011100000000001",--11259
"001111001100000010000000000000000010",--11260
"010110010001000001110000000000000010",--11261
"001111010000000001110000000000000011",--11262
"011110001111000000000000000000010011",--11263
"001111010000000001100000000000000100",--11264
"111110001100010001010010100000000000",--11265
"001111010000000001100000000000000101",--11266
"111110001010001001100010100000000000",--11267
"001111001110000001100000000000000000",--11268
"111110001010001001100011000000000000",--11269
"111110001100000000110001100000000001",--11270
"001111001100000001100000000000000000",--11271
"010110001101000000110000000000110110",--11272
"001111001110000000110000000000000001",--11273
"111110001010001000110001100000000000",--11274
"111110000110000001000001100000000001",--11275
"001111001100000001000000000000000001",--11276
"010110001001000000110000000000110001",--11277
"001111010000000000110000000000000101",--11278
"010010000111000000000000000000101111",--11279
"001011000000000001010000000100101111",--11280
"101001000000000001100000000000000011",--11281
"000101000000000000000010110001001010",--11282
"001011000000000001100000000100101111",--11283
"101001000000000001100000000000000010",--11284
"000101000000000000000010110001001010",--11285
"001011000000000001100000000100101111",--11286
"101001000000000001100000000000000001",--11287
"000101000000000000000010110001001010",--11288
"011111010011000000100000000000000111",--11289
"001111010000000000110000000000000000",--11290
"011010000111000000000000000000100011",--11291
"001111001110000001000000000000000011",--11292
"111110000110001001000001100000000000",--11293
"001011000000000000110000000100101111",--11294
"101001000000000001100000000000000001",--11295
"000101000000000000000010110001001010",--11296
"001111010000000001100000000000000000",--11297
"010010001101000000000000000000011100",--11298
"001111010000000001110000000000000001",--11299
"111110001110001000110001100000000000",--11300
"001111010000000001110000000000000010",--11301
"111110001110001001000010000000000000",--11302
"111110000110000001000001100000000000",--11303
"001111010000000001000000000000000011",--11304
"111110001000001001010010000000000000",--11305
"111110000110000001000001100000000000",--11306
"001111001110000001000000000000000011",--11307
"111110000110001000110010100000000000",--11308
"111110001100001001000010000000000000",--11309
"111110001010010001000010000000000000",--11310
"010110001001000000000000000000001111",--11311
"001101001100000001100000000000000110",--11312
"011100001101000000000000000000000110",--11313
"111110001000100000000010000000000000",--11314
"111110000110010001000001100000000000",--11315
"001111010000000001000000000000000100",--11316
"111110000110001001000001100000000000",--11317
"001011000000000000110000000100101111",--11318
"000101000000000000000010110000111101",--11319
"111110001000100000000010000000000000",--11320
"111110000110000001000001100000000000",--11321
"001111010000000001000000000000000100",--11322
"111110000110001001000001100000000000",--11323
"001011000000000000110000000100101111",--11324
"101001000000000001100000000000000001",--11325
"000101000000000000000010110001001010",--11326
"001101001010000001010000000101101101",--11327
"001101001010000001010000000000000110",--11328
"010000001011000000000000000011100100",--11329
"101000001001111000000001000000000000",--11330
"101001000000000000010000000000000001",--11331
"001001111100000111111111111111111101",--11332
"101001111100010111100000000000000100",--11333
"000111000000000000000010011110011001",--11334
"101001111100000111100000000000000100",--11335
"001101111100000111111111111111111101",--11336
"000101000000000000000010110100100110",--11337
"001111000000000000110000000100101111",--11338
"001001111100000001001111111111111101",--11339
"010110000111000000000000000011010001",--11340
"001111000000000001000000000100101101",--11341
"010110001001000000110000000011001111",--11342
"001101000110000001110000000000000000",--11343
"101111001001110001000011110000100011",--11344
"101111001001100001001101011100001010",--11345
"111110000110000001000001100000000000",--11346
"001111001110000001000000000000000000",--11347
"111110001000001000110010000000000000",--11348
"001111000000000001010000000100010010",--11349
"111110001000000001010010000000000000",--11350
"001111001110000001010000000000000001",--11351
"111110001010001000110010100000000000",--11352
"001111000000000001100000000100010011",--11353
"111110001010000001100010100000000000",--11354
"001111001110000001100000000000000010",--11355
"111110001100001000110011000000000000",--11356
"001111000000000001110000000100010100",--11357
"111110001100000001110011000000000000",--11358
"001101001000000001110000000000000000",--11359
"001001111100000001101111111111111100",--11360
"001001111100000001011111111111111011",--11361
"001011111100000001101111111111111010",--11362
"001011111100000001011111111111111001",--11363
"001011111100000001001111111111111000",--11364
"001011111100000000111111111111110111",--11365
"010011001111000000000000000010101011",--11366
"001101001110000001110000000101101101",--11367
"001101001110000010000000000000000101",--11368
"001111010000000001110000000000000000",--11369
"111110001000010001110011100000000000",--11370
"001111010000000010000000000000000001",--11371
"111110001010010010000100000000000000",--11372
"001111010000000010010000000000000010",--11373
"111110001100010010010100100000000000",--11374
"001101001110000010000000000000000001",--11375
"011111010001000000010000000000010000",--11376
"101110001111111000000011100000000001",--11377
"001101001110000010000000000000000100",--11378
"001111010000000010100000000000000000",--11379
"010110010101000001110000000000001001",--11380
"101110010001111000000011100000000001",--11381
"001111010000000010000000000000000001",--11382
"010110010001000001110000000000000110",--11383
"101110010011111000000011100000000001",--11384
"001111010000000010000000000000000010",--11385
"010110010001000001110000000000000011",--11386
"001101001110000001110000000000000110",--11387
"011100001111000000000000000010100001",--11388
"000101000000000000000010110010110110",--11389
"001101001110000001110000000000000110",--11390
"011100001111000000000000000000110110",--11391
"000101000000000000000010110100011110",--11392
"011111010001000000100000000000001111",--11393
"001101001110000010000000000000000100",--11394
"001111010000000010100000000000000000",--11395
"111110010100001001110011100000000000",--11396
"001111010000000010100000000000000001",--11397
"111110010100001010000100000000000000",--11398
"111110001110000010000011100000000000",--11399
"001111010000000010000000000000000010",--11400
"111110010000001010010100000000000000",--11401
"111110001110000010000011100000000000",--11402
"001101001110000001110000000000000110",--11403
"011010001111000000000000000000000010",--11404
"011111001111000000010000000000101000",--11405
"000101000000000000000010110100011110",--11406
"011100001111000000000000000000100110",--11407
"000101000000000000000010110100011110",--11408
"111110001110001001110101000000000000",--11409
"001101001110000010010000000000000100",--11410
"001111010010000010110000000000000000",--11411
"111110010100001010110101000000000000",--11412
"111110010000001010000101100000000000",--11413
"001111010010000011000000000000000001",--11414
"111110010110001011000101100000000000",--11415
"111110010100000010110101000000000000",--11416
"111110010010001010010101100000000000",--11417
"001111010010000011000000000000000010",--11418
"111110010110001011000101100000000000",--11419
"111110010100000010110101000000000000",--11420
"001101001110000010010000000000000011",--11421
"011100010011000000000000000000000011",--11422
"101110010101111000000011100000000000",--11423
"011111010001000000110000000000010000",--11424
"000101000000000000000010110010110000",--11425
"111110010000001010010101100000000000",--11426
"001101001110000010010000000000001001",--11427
"001111010010000011000000000000000000",--11428
"111110010110001011000101100000000000",--11429
"111110010100000010110101000000000000",--11430
"111110010010001001110100100000000000",--11431
"001111010010000010110000000000000001",--11432
"111110010010001010110100100000000000",--11433
"111110010100000010010100100000000000",--11434
"111110001110001010000011100000000000",--11435
"001111010010000010000000000000000010",--11436
"111110001110001010000011100000000000",--11437
"111110010010000001110011100000000000",--11438
"011111010001000000110000000000000001",--11439
"111110001110010000010011100000000000",--11440
"001101001110000001110000000000000110",--11441
"011010001111000000000000000000000010",--11442
"011111001111000000010000000000000010",--11443
"000101000000000000000010110100011110",--11444
"010000001111000000000000000001101000",--11445
"001101001000000001110000000000000001",--11446
"010011001111000000000000000001011010",--11447
"001101001110000001110000000101101101",--11448
"001101001110000010000000000000000101",--11449
"001111010000000001110000000000000000",--11450
"111110001000010001110011100000000000",--11451
"001111010000000010000000000000000001",--11452
"111110001010010010000100000000000000",--11453
"001111010000000010010000000000000010",--11454
"111110001100010010010100100000000000",--11455
"001101001110000010000000000000000001",--11456
"011111010001000000010000000000010000",--11457
"101110001111111000000011100000000001",--11458
"001101001110000010000000000000000100",--11459
"001111010000000010100000000000000000",--11460
"010110010101000001110000000000001001",--11461
"101110010001111000000011100000000001",--11462
"001111010000000010000000000000000001",--11463
"010110010001000001110000000000000110",--11464
"101110010011111000000011100000000001",--11465
"001111010000000010000000000000000010",--11466
"010110010001000001110000000000000011",--11467
"001101001110000001110000000000000110",--11468
"011100001111000000000000000001010000",--11469
"000101000000000000000010110100000111",--11470
"001101001110000001110000000000000110",--11471
"011100001111000000000000000000110110",--11472
"000101000000000000000010110100011110",--11473
"011111010001000000100000000000001111",--11474
"001101001110000010000000000000000100",--11475
"001111010000000010100000000000000000",--11476
"111110010100001001110011100000000000",--11477
"001111010000000010100000000000000001",--11478
"111110010100001010000100000000000000",--11479
"111110001110000010000011100000000000",--11480
"001111010000000010000000000000000010",--11481
"111110010000001010010100000000000000",--11482
"111110001110000010000011100000000000",--11483
"001101001110000001110000000000000110",--11484
"011010001111000000000000000000000010",--11485
"011111001111000000010000000000101000",--11486
"000101000000000000000010110100011110",--11487
"011100001111000000000000000000100110",--11488
"000101000000000000000010110100011110",--11489
"111110001110001001110101000000000000",--11490
"001101001110000010010000000000000100",--11491
"001111010010000010110000000000000000",--11492
"111110010100001010110101000000000000",--11493
"111110010000001010000101100000000000",--11494
"001111010010000011000000000000000001",--11495
"111110010110001011000101100000000000",--11496
"111110010100000010110101000000000000",--11497
"111110010010001010010101100000000000",--11498
"001111010010000011000000000000000010",--11499
"111110010110001011000101100000000000",--11500
"111110010100000010110101000000000000",--11501
"001101001110000010010000000000000011",--11502
"011100010011000000000000000000000011",--11503
"101110010101111000000011100000000000",--11504
"011111010001000000110000000000010000",--11505
"000101000000000000000010110100000001",--11506
"111110010000001010010101100000000000",--11507
"001101001110000010010000000000001001",--11508
"001111010010000011000000000000000000",--11509
"111110010110001011000101100000000000",--11510
"111110010100000010110101000000000000",--11511
"111110010010001001110100100000000000",--11512
"001111010010000010110000000000000001",--11513
"111110010010001010110100100000000000",--11514
"111110010100000010010100100000000000",--11515
"111110001110001010000011100000000000",--11516
"001111010010000010000000000000000010",--11517
"111110001110001010000011100000000000",--11518
"111110010010000001110011100000000000",--11519
"011111010001000000110000000000000001",--11520
"111110001110010000010011100000000000",--11521
"001101001110000001110000000000000110",--11522
"011010001111000000000000000000000010",--11523
"011111001111000000010000000000000010",--11524
"000101000000000000000010110100011110",--11525
"010000001111000000000000000000010111",--11526
"101000001001111000000001000000000000",--11527
"101001000000000000010000000000000010",--11528
"101110001001111000000001100000000000",--11529
"101110001011111000000010000000000000",--11530
"101110001101111000000010100000000000",--11531
"001001111100000111111111111111110110",--11532
"101001111100010111100000000000001011",--11533
"000111000000000000000000011110001000",--11534
"101001111100000111100000000000001011",--11535
"001101111100000111111111111111110110",--11536
"010000000011000000000000000000001100",--11537
"001111111100000000111111111111110111",--11538
"001011000000000000110000000100101101",--11539
"001111111100000000111111111111111000",--11540
"001011000000000000110000000100101010",--11541
"001111111100000000111111111111111001",--11542
"001011000000000000110000000100101011",--11543
"001111111100000000111111111111111010",--11544
"001011000000000000110000000100101100",--11545
"001101111100000000011111111111111011",--11546
"001001000000000000010000000100101001",--11547
"001101111100000000011111111111111100",--11548
"001001000000000000010000000100101110",--11549
"101001000000000000010000000000000001",--11550
"001101111100000000101111111111111101",--11551
"001101111100000000110000000000000000",--11552
"001001111100000111111111111111111100",--11553
"101001111100010111100000000000000101",--11554
"000111000000000000000010011110011001",--11555
"101001111100000111100000000000000101",--11556
"001101111100000111111111111111111100",--11557
"001101111100000000011111111111111110",--11558
"101001000010000000010000000000000001",--11559
"001101111100000000111111111111111111",--11560
"001100000110000000010001000000000000",--11561
"010011000100000000001111100000000000",--11562
"001101000100000000100000000100110001",--11563
"001101111100000000110000000000000000",--11564
"001001111100000000011111111111111101",--11565
"101000000001111000000000100000000000",--11566
"001001111100000111111111111111111100",--11567
"101001111100010111100000000000000101",--11568
"000111000000000000000010011110011001",--11569
"101001111100000111100000000000000101",--11570
"001101111100000111111111111111111100",--11571
"001101111100000000011111111111111101",--11572
"101001000010000000010000000000000001",--11573
"001101111100000000111111111111111111",--11574
"001100000110000000010001000000000000",--11575
"010011000100000000001111100000000000",--11576
"001101000100000000100000000100110001",--11577
"001101000100000001000000000000000000",--11578
"001001111100000000011111111111111100",--11579
"010011001001000000000000000010101111",--11580
"001101001000000001010000000101101101",--11581
"001101001010000001100000000000001010",--11582
"001111001100000000110000000000000000",--11583
"001111001100000001000000000000000001",--11584
"001111001100000001010000000000000010",--11585
"001101111100000001110000000000000000",--11586
"001101001110000010000000000000000001",--11587
"001100010000000001000100000000000000",--11588
"001101001010000010010000000000000001",--11589
"011111010011000000010000000000111011",--11590
"001101001110000001100000000000000000",--11591
"001111010000000001100000000000000000",--11592
"111110001100010000110011000000000000",--11593
"001111010000000001110000000000000001",--11594
"111110001100001001110011000000000000",--11595
"001111001100000001110000000000000001",--11596
"111110001100001001110011100000000000",--11597
"111110001110000001000011100000000001",--11598
"001101001010000001010000000000000100",--11599
"001111001010000010000000000000000001",--11600
"010110010001000001110000000000000111",--11601
"001111001100000001110000000000000010",--11602
"111110001100001001110011100000000000",--11603
"111110001110000001010011100000000001",--11604
"001111001010000010000000000000000010",--11605
"010110010001000001110000000000000010",--11606
"001111010000000001110000000000000001",--11607
"011110001111000000000000000000100110",--11608
"001111010000000001100000000000000010",--11609
"111110001100010001000011000000000000",--11610
"001111010000000001110000000000000011",--11611
"111110001100001001110011000000000000",--11612
"001111001100000001110000000000000000",--11613
"111110001100001001110011100000000000",--11614
"111110001110000000110011100000000001",--11615
"001111001010000010000000000000000000",--11616
"010110010001000001110000000000000111",--11617
"001111001100000001110000000000000010",--11618
"111110001100001001110011100000000000",--11619
"111110001110000001010011100000000001",--11620
"001111001010000010000000000000000010",--11621
"010110010001000001110000000000000010",--11622
"001111010000000001110000000000000011",--11623
"011110001111000000000000000000010011",--11624
"001111010000000001100000000000000100",--11625
"111110001100010001010010100000000000",--11626
"001111010000000001100000000000000101",--11627
"111110001010001001100010100000000000",--11628
"001111001100000001100000000000000000",--11629
"111110001010001001100011000000000000",--11630
"111110001100000000110001100000000001",--11631
"001111001010000001100000000000000000",--11632
"010110001101000000110000000000110110",--11633
"001111001100000000110000000000000001",--11634
"111110001010001000110001100000000000",--11635
"111110000110000001000001100000000001",--11636
"001111001010000001000000000000000001",--11637
"010110001001000000110000000000110001",--11638
"001111010000000000110000000000000101",--11639
"010010000111000000000000000000101111",--11640
"001011000000000001010000000100101111",--11641
"101001000000000001010000000000000011",--11642
"000101000000000000000010110110110011",--11643
"001011000000000001100000000100101111",--11644
"101001000000000001010000000000000010",--11645
"000101000000000000000010110110110011",--11646
"001011000000000001100000000100101111",--11647
"101001000000000001010000000000000001",--11648
"000101000000000000000010110110110011",--11649
"011111010011000000100000000000000111",--11650
"001111010000000000110000000000000000",--11651
"011010000111000000000000000000100011",--11652
"001111001100000001000000000000000011",--11653
"111110000110001001000001100000000000",--11654
"001011000000000000110000000100101111",--11655
"101001000000000001010000000000000001",--11656
"000101000000000000000010110110110011",--11657
"001111010000000001100000000000000000",--11658
"010010001101000000000000000000011100",--11659
"001111010000000001110000000000000001",--11660
"111110001110001000110001100000000000",--11661
"001111010000000001110000000000000010",--11662
"111110001110001001000010000000000000",--11663
"111110000110000001000001100000000000",--11664
"001111010000000001000000000000000011",--11665
"111110001000001001010010000000000000",--11666
"111110000110000001000001100000000000",--11667
"001111001100000001000000000000000011",--11668
"111110000110001000110010100000000000",--11669
"111110001100001001000010000000000000",--11670
"111110001010010001000010000000000000",--11671
"010110001001000000000000000000001111",--11672
"001101001010000001010000000000000110",--11673
"011100001011000000000000000000000110",--11674
"111110001000100000000010000000000000",--11675
"111110000110010001000001100000000000",--11676
"001111010000000001000000000000000100",--11677
"111110000110001001000001100000000000",--11678
"001011000000000000110000000100101111",--11679
"000101000000000000000010110110100110",--11680
"111110001000100000000010000000000000",--11681
"111110000110000001000001100000000000",--11682
"001111010000000001000000000000000100",--11683
"111110000110001001000001100000000000",--11684
"001011000000000000110000000100101111",--11685
"101001000000000001010000000000000001",--11686
"000101000000000000000010110110110011",--11687
"001101001000000001000000000101101101",--11688
"001101001000000001000000000000000110",--11689
"010000001001000000000000000001000001",--11690
"101000001111111000000001100000000000",--11691
"101001000000000000010000000000000001",--11692
"001001111100000111111111111111111011",--11693
"101001111100010111100000000000000110",--11694
"000111000000000000000010011110011001",--11695
"101001111100000111100000000000000110",--11696
"001101111100000111111111111111111011",--11697
"000101000000000000000010110111101100",--11698
"001111000000000000110000000100101111",--11699
"001001111100000000101111111111111011",--11700
"010110000111000000000000000000101110",--11701
"001111000000000001000000000100101101",--11702
"010110001001000000110000000000101100",--11703
"001101001110000001100000000000000000",--11704
"101111001001110001000011110000100011",--11705
"101111001001100001001101011100001010",--11706
"111110000110000001000001100000000000",--11707
"001111001100000001000000000000000000",--11708
"111110001000001000110010000000000000",--11709
"001111000000000001010000000100010010",--11710
"111110001000000001010010000000000000",--11711
"001111001100000001010000000000000001",--11712
"111110001010001000110010100000000000",--11713
"001111000000000001100000000100010011",--11714
"111110001010000001100010100000000000",--11715
"001111001100000001100000000000000010",--11716
"111110001100001000110011000000000000",--11717
"001111000000000001110000000100010100",--11718
"111110001100000001110011000000000000",--11719
"001001111100000001011111111111111010",--11720
"001001111100000001001111111111111001",--11721
"001011111100000001101111111111111000",--11722
"001011111100000001011111111111110111",--11723
"001011111100000001001111111111110110",--11724
"001011111100000000111111111111110101",--11725
"101000000001111000000000100000000000",--11726
"101110001001111000000001100000000000",--11727
"101110001011111000000010000000000000",--11728
"101110001101111000000010100000000000",--11729
"001001111100000111111111111111110100",--11730
"101001111100010111100000000000001101",--11731
"000111000000000000000000011110001000",--11732
"101001111100000111100000000000001101",--11733
"001101111100000111111111111111110100",--11734
"010000000011000000000000000000001100",--11735
"001111111100000000111111111111110101",--11736
"001011000000000000110000000100101101",--11737
"001111111100000000111111111111110110",--11738
"001011000000000000110000000100101010",--11739
"001111111100000000111111111111110111",--11740
"001011000000000000110000000100101011",--11741
"001111111100000000111111111111111000",--11742
"001011000000000000110000000100101100",--11743
"001101111100000000011111111111111001",--11744
"001001000000000000010000000100101001",--11745
"001101111100000000011111111111111010",--11746
"001001000000000000010000000100101110",--11747
"101001000000000000010000000000000001",--11748
"001101111100000000101111111111111011",--11749
"001101111100000000110000000000000000",--11750
"001001111100000111111111111111111010",--11751
"101001111100010111100000000000000111",--11752
"000111000000000000000010011110011001",--11753
"101001111100000111100000000000000111",--11754
"001101111100000111111111111111111010",--11755
"001101111100000000011111111111111100",--11756
"101001000010000000010000000000000001",--11757
"001101111100000000111111111111111111",--11758
"001100000110000000010001000000000000",--11759
"010011000100000000001111100000000000",--11760
"001101000100000000100000000100110001",--11761
"001101111100000000110000000000000000",--11762
"001001111100000000011111111111111011",--11763
"101000000001111000000000100000000000",--11764
"001001111100000111111111111111111010",--11765
"101001111100010111100000000000000111",--11766
"000111000000000000000010011110011001",--11767
"101001111100000111100000000000000111",--11768
"001101111100000111111111111111111010",--11769
"001101111100000000011111111111111011",--11770
"101001000010000000010000000000000001",--11771
"001101111100000000101111111111111111",--11772
"001101111100000000110000000000000000",--11773
"000101000000000000000010101111001101",--11774
"001100000100000000010010000000000000",--11775
"001101001000000001010000000000000000",--11776
"010011001010000000001111100000000000",--11777
"001001111100000000110000000000000000",--11778
"001001111100000000101111111111111111",--11779
"001001111100000000011111111111111110",--11780
"011111001011011000110000000011010001",--11781
"001101001000000001010000000000000001",--11782
"010011001011000000000000001000001000",--11783
"001101001010000000100000000100110001",--11784
"001001111100000001001111111111111101",--11785
"101000000001111000000000100000000000",--11786
"001001111100000111111111111111111100",--11787
"101001111100010111100000000000000101",--11788
"000111000000000000000010011110011001",--11789
"101001111100000111100000000000000101",--11790
"001101111100000111111111111111111100",--11791
"001101111100000000011111111111111101",--11792
"001101000010000000100000000000000010",--11793
"010011000101000000000000000111111101",--11794
"001101000100000000100000000100110001",--11795
"001101000100000000110000000000000000",--11796
"010011000111000000000000000010101111",--11797
"001101000110000001000000000101101101",--11798
"001101001000000001010000000000001010",--11799
"001111001010000000110000000000000000",--11800
"001111001010000001000000000000000001",--11801
"001111001010000001010000000000000010",--11802
"001101111100000001100000000000000000",--11803
"001101001100000001110000000000000001",--11804
"001100001110000000110011100000000000",--11805
"001101001000000010000000000000000001",--11806
"011111010001000000010000000000111011",--11807
"001101001100000001010000000000000000",--11808
"001111001110000001100000000000000000",--11809
"111110001100010000110011000000000000",--11810
"001111001110000001110000000000000001",--11811
"111110001100001001110011000000000000",--11812
"001111001010000001110000000000000001",--11813
"111110001100001001110011100000000000",--11814
"111110001110000001000011100000000001",--11815
"001101001000000001000000000000000100",--11816
"001111001000000010000000000000000001",--11817
"010110010001000001110000000000000111",--11818
"001111001010000001110000000000000010",--11819
"111110001100001001110011100000000000",--11820
"111110001110000001010011100000000001",--11821
"001111001000000010000000000000000010",--11822
"010110010001000001110000000000000010",--11823
"001111001110000001110000000000000001",--11824
"011110001111000000000000000000100110",--11825
"001111001110000001100000000000000010",--11826
"111110001100010001000011000000000000",--11827
"001111001110000001110000000000000011",--11828
"111110001100001001110011000000000000",--11829
"001111001010000001110000000000000000",--11830
"111110001100001001110011100000000000",--11831
"111110001110000000110011100000000001",--11832
"001111001000000010000000000000000000",--11833
"010110010001000001110000000000000111",--11834
"001111001010000001110000000000000010",--11835
"111110001100001001110011100000000000",--11836
"111110001110000001010011100000000001",--11837
"001111001000000010000000000000000010",--11838
"010110010001000001110000000000000010",--11839
"001111001110000001110000000000000011",--11840
"011110001111000000000000000000010011",--11841
"001111001110000001100000000000000100",--11842
"111110001100010001010010100000000000",--11843
"001111001110000001100000000000000101",--11844
"111110001010001001100010100000000000",--11845
"001111001010000001100000000000000000",--11846
"111110001010001001100011000000000000",--11847
"111110001100000000110001100000000001",--11848
"001111001000000001100000000000000000",--11849
"010110001101000000110000000000110110",--11850
"001111001010000000110000000000000001",--11851
"111110001010001000110001100000000000",--11852
"111110000110000001000001100000000001",--11853
"001111001000000001000000000000000001",--11854
"010110001001000000110000000000110001",--11855
"001111001110000000110000000000000101",--11856
"010010000111000000000000000000101111",--11857
"001011000000000001010000000100101111",--11858
"101001000000000001000000000000000011",--11859
"000101000000000000000010111010001100",--11860
"001011000000000001100000000100101111",--11861
"101001000000000001000000000000000010",--11862
"000101000000000000000010111010001100",--11863
"001011000000000001100000000100101111",--11864
"101001000000000001000000000000000001",--11865
"000101000000000000000010111010001100",--11866
"011111010001000000100000000000000111",--11867
"001111001110000000110000000000000000",--11868
"011010000111000000000000000000100011",--11869
"001111001010000001000000000000000011",--11870
"111110000110001001000001100000000000",--11871
"001011000000000000110000000100101111",--11872
"101001000000000001000000000000000001",--11873
"000101000000000000000010111010001100",--11874
"001111001110000001100000000000000000",--11875
"010010001101000000000000000000011100",--11876
"001111001110000001110000000000000001",--11877
"111110001110001000110001100000000000",--11878
"001111001110000001110000000000000010",--11879
"111110001110001001000010000000000000",--11880
"111110000110000001000001100000000000",--11881
"001111001110000001000000000000000011",--11882
"111110001000001001010010000000000000",--11883
"111110000110000001000001100000000000",--11884
"001111001010000001000000000000000011",--11885
"111110000110001000110010100000000000",--11886
"111110001100001001000010000000000000",--11887
"111110001010010001000010000000000000",--11888
"010110001001000000000000000000001111",--11889
"001101001000000001000000000000000110",--11890
"011100001001000000000000000000000110",--11891
"111110001000100000000010000000000000",--11892
"111110000110010001000001100000000000",--11893
"001111001110000001000000000000000100",--11894
"111110000110001001000001100000000000",--11895
"001011000000000000110000000100101111",--11896
"000101000000000000000010111001111111",--11897
"111110001000100000000010000000000000",--11898
"111110000110000001000001100000000000",--11899
"001111001110000001000000000000000100",--11900
"111110000110001001000001100000000000",--11901
"001011000000000000110000000100101111",--11902
"101001000000000001000000000000000001",--11903
"000101000000000000000010111010001100",--11904
"001101000110000000110000000101101101",--11905
"001101000110000000110000000000000110",--11906
"010000000111000000000000000001000001",--11907
"101001000000000000010000000000000001",--11908
"101000001101111000000001100000000000",--11909
"001001111100000111111111111111111100",--11910
"101001111100010111100000000000000101",--11911
"000111000000000000000010011110011001",--11912
"101001111100000111100000000000000101",--11913
"001101111100000111111111111111111100",--11914
"000101000000000000000010111011000101",--11915
"001111000000000000110000000100101111",--11916
"001001111100000000101111111111111100",--11917
"010110000111000000000000000000101110",--11918
"001111000000000001000000000100101101",--11919
"010110001001000000110000000000101100",--11920
"001101001100000001010000000000000000",--11921
"101111001001110001000011110000100011",--11922
"101111001001100001001101011100001010",--11923
"111110000110000001000001100000000000",--11924
"001111001010000001000000000000000000",--11925
"111110001000001000110010000000000000",--11926
"001111000000000001010000000100010010",--11927
"111110001000000001010010000000000000",--11928
"001111001010000001010000000000000001",--11929
"111110001010001000110010100000000000",--11930
"001111000000000001100000000100010011",--11931
"111110001010000001100010100000000000",--11932
"001111001010000001100000000000000010",--11933
"111110001100001000110011000000000000",--11934
"001111000000000001110000000100010100",--11935
"111110001100000001110011000000000000",--11936
"001001111100000001001111111111111011",--11937
"001001111100000000111111111111111010",--11938
"001011111100000001101111111111111001",--11939
"001011111100000001011111111111111000",--11940
"001011111100000001001111111111110111",--11941
"001011111100000000111111111111110110",--11942
"101000000001111000000000100000000000",--11943
"101110001001111000000001100000000000",--11944
"101110001011111000000010000000000000",--11945
"101110001101111000000010100000000000",--11946
"001001111100000111111111111111110101",--11947
"101001111100010111100000000000001100",--11948
"000111000000000000000000011110001000",--11949
"101001111100000111100000000000001100",--11950
"001101111100000111111111111111110101",--11951
"010000000011000000000000000000001100",--11952
"001111111100000000111111111111110110",--11953
"001011000000000000110000000100101101",--11954
"001111111100000000111111111111110111",--11955
"001011000000000000110000000100101010",--11956
"001111111100000000111111111111111000",--11957
"001011000000000000110000000100101011",--11958
"001111111100000000111111111111111001",--11959
"001011000000000000110000000100101100",--11960
"001101111100000000011111111111111010",--11961
"001001000000000000010000000100101001",--11962
"001101111100000000011111111111111011",--11963
"001001000000000000010000000100101110",--11964
"101001000000000000010000000000000001",--11965
"001101111100000000101111111111111100",--11966
"001101111100000000110000000000000000",--11967
"001001111100000111111111111111111011",--11968
"101001111100010111100000000000000110",--11969
"000111000000000000000010011110011001",--11970
"101001111100000111100000000000000110",--11971
"001101111100000111111111111111111011",--11972
"001101111100000000011111111111111101",--11973
"001101000010000000100000000000000011",--11974
"010011000101000000000000000101001000",--11975
"001101000100000000100000000100110001",--11976
"001101111100000000110000000000000000",--11977
"101000000001111000000000100000000000",--11978
"001001111100000111111111111111111100",--11979
"101001111100010111100000000000000101",--11980
"000111000000000000000010011110011001",--11981
"101001111100000111100000000000000101",--11982
"101001000000000000010000000000000100",--11983
"001101111100000000101111111111111101",--11984
"001101111100000000110000000000000000",--11985
"101001111100010111100000000000000101",--11986
"000111000000000000000010101111001101",--11987
"101001111100000111100000000000000101",--11988
"001101111100000111111111111111111100",--11989
"000101000000000000000011000000010000",--11990
"001101001010000001100000000101101101",--11991
"001101001100000001110000000000001010",--11992
"001111001110000000110000000000000000",--11993
"001111001110000001000000000000000001",--11994
"001111001110000001010000000000000010",--11995
"001101000110000010000000000000000001",--11996
"001100010000000001010010100000000000",--11997
"001101001100000010010000000000000001",--11998
"011111010011000000010000000000111000",--11999
"001101000110000001110000000000000000",--12000
"001111001010000001100000000000000000",--12001
"111110001100010000110011000000000000",--12002
"001111001010000001110000000000000001",--12003
"111110001100001001110011000000000000",--12004
"001111001110000001110000000000000001",--12005
"111110001100001001110011100000000000",--12006
"111110001110000001000011100000000001",--12007
"001101001100000001100000000000000100",--12008
"001111001100000010000000000000000001",--12009
"010110010001000001110000000000000111",--12010
"001111001110000001110000000000000010",--12011
"111110001100001001110011100000000000",--12012
"111110001110000001010011100000000001",--12013
"001111001100000010000000000000000010",--12014
"010110010001000001110000000000000010",--12015
"001111001010000001110000000000000001",--12016
"011110001111000000000000000000100100",--12017
"001111001010000001100000000000000010",--12018
"111110001100010001000011000000000000",--12019
"001111001010000001110000000000000011",--12020
"111110001100001001110011000000000000",--12021
"001111001110000001110000000000000000",--12022
"111110001100001001110011100000000000",--12023
"111110001110000000110011100000000001",--12024
"001111001100000010000000000000000000",--12025
"010110010001000001110000000000000111",--12026
"001111001110000001110000000000000010",--12027
"111110001100001001110011100000000000",--12028
"111110001110000001010011100000000001",--12029
"001111001100000010000000000000000010",--12030
"010110010001000001110000000000000010",--12031
"001111001010000001110000000000000011",--12032
"011110001111000000000000000000010010",--12033
"001111001010000001100000000000000100",--12034
"111110001100010001010010100000000000",--12035
"001111001010000001100000000000000101",--12036
"111110001010001001100010100000000000",--12037
"001111001110000001100000000000000000",--12038
"111110001010001001100011000000000000",--12039
"111110001100000000110001100000000001",--12040
"001111001100000001100000000000000000",--12041
"010110001101000000110000000100000101",--12042
"001111001110000000110000000000000001",--12043
"111110001010001000110001100000000000",--12044
"111110000110000001000001100000000001",--12045
"001111001100000001000000000000000001",--12046
"010110001001000000110000000100000000",--12047
"001111001010000000110000000000000101",--12048
"010010000111000000000000000011111110",--12049
"001011000000000001010000000100101111",--12050
"000101000000000000000010111100111011",--12051
"001011000000000001100000000100101111",--12052
"000101000000000000000010111100111011",--12053
"001011000000000001100000000100101111",--12054
"000101000000000000000010111100111011",--12055
"011111010011000000100000000000000110",--12056
"001111001010000000110000000000000000",--12057
"011010000111000000000000000011110101",--12058
"001111001110000001000000000000000011",--12059
"111110000110001001000001100000000000",--12060
"001011000000000000110000000100101111",--12061
"000101000000000000000010111100111011",--12062
"001111001010000001100000000000000000",--12063
"010010001101000000000000000011101111",--12064
"001111001010000001110000000000000001",--12065
"111110001110001000110001100000000000",--12066
"001111001010000001110000000000000010",--12067
"111110001110001001000010000000000000",--12068
"111110000110000001000001100000000000",--12069
"001111001010000001000000000000000011",--12070
"111110001000001001010010000000000000",--12071
"111110000110000001000001100000000000",--12072
"001111001110000001000000000000000011",--12073
"111110000110001000110010100000000000",--12074
"111110001100001001000010000000000000",--12075
"111110001010010001000010000000000000",--12076
"010110001001000000000000000011100010",--12077
"001101001100000001100000000000000110",--12078
"011100001101000000000000000000000110",--12079
"111110001000100000000010000000000000",--12080
"111110000110010001000001100000000000",--12081
"001111001010000001000000000000000100",--12082
"111110000110001001000001100000000000",--12083
"001011000000000000110000000100101111",--12084
"000101000000000000000010111100111011",--12085
"111110001000100000000010000000000000",--12086
"111110000110000001000001100000000000",--12087
"001111001010000001000000000000000100",--12088
"111110000110001001000001100000000000",--12089
"001011000000000000110000000100101111",--12090
"001111000000000000110000000100101111",--12091
"001111000000000001000000000100101101",--12092
"010110001001000000110000000011010010",--12093
"001101001000000001010000000000000001",--12094
"010011001011000000000000000011010000",--12095
"001101001010000000100000000100110001",--12096
"001001111100000010001111111111111101",--12097
"001001111100000001001111111111111100",--12098
"101000000001111000000000100000000000",--12099
"001001111100000111111111111111111011",--12100
"101001111100010111100000000000000110",--12101
"000111000000000000000010011110011001",--12102
"101001111100000111100000000000000110",--12103
"001101111100000111111111111111111011",--12104
"001101111100000000011111111111111100",--12105
"001101000010000000100000000000000010",--12106
"010011000101000000000000000011000100",--12107
"001101000100000000100000000100110001",--12108
"001101000100000000110000000000000000",--12109
"010011000111000000000000000010110000",--12110
"001101000110000001000000000101101101",--12111
"001101001000000001010000000000001010",--12112
"001111001010000000110000000000000000",--12113
"001111001010000001000000000000000001",--12114
"001111001010000001010000000000000010",--12115
"001101111100000001111111111111111101",--12116
"001100001110000000110011000000000000",--12117
"001101001000000001110000000000000001",--12118
"011111001111000000010000000000111100",--12119
"001101111100000001010000000000000000",--12120
"001101001010000001110000000000000000",--12121
"001111001100000001100000000000000000",--12122
"111110001100010000110011000000000000",--12123
"001111001100000001110000000000000001",--12124
"111110001100001001110011000000000000",--12125
"001111001110000001110000000000000001",--12126
"111110001100001001110011100000000000",--12127
"111110001110000001000011100000000001",--12128
"001101001000000001000000000000000100",--12129
"001111001000000010000000000000000001",--12130
"010110010001000001110000000000000111",--12131
"001111001110000001110000000000000010",--12132
"111110001100001001110011100000000000",--12133
"111110001110000001010011100000000001",--12134
"001111001000000010000000000000000010",--12135
"010110010001000001110000000000000010",--12136
"001111001100000001110000000000000001",--12137
"011110001111000000000000000000100110",--12138
"001111001100000001100000000000000010",--12139
"111110001100010001000011000000000000",--12140
"001111001100000001110000000000000011",--12141
"111110001100001001110011000000000000",--12142
"001111001110000001110000000000000000",--12143
"111110001100001001110011100000000000",--12144
"111110001110000000110011100000000001",--12145
"001111001000000010000000000000000000",--12146
"010110010001000001110000000000000111",--12147
"001111001110000001110000000000000010",--12148
"111110001100001001110011100000000000",--12149
"111110001110000001010011100000000001",--12150
"001111001000000010000000000000000010",--12151
"010110010001000001110000000000000010",--12152
"001111001100000001110000000000000011",--12153
"011110001111000000000000000000010011",--12154
"001111001100000001100000000000000100",--12155
"111110001100010001010010100000000000",--12156
"001111001100000001100000000000000101",--12157
"111110001010001001100010100000000000",--12158
"001111001110000001100000000000000000",--12159
"111110001010001001100011000000000000",--12160
"111110001100000000110001100000000001",--12161
"001111001000000001100000000000000000",--12162
"010110001101000000110000000000110110",--12163
"001111001110000000110000000000000001",--12164
"111110001010001000110001100000000000",--12165
"111110000110000001000001100000000001",--12166
"001111001000000001000000000000000001",--12167
"010110001001000000110000000000110001",--12168
"001111001100000000110000000000000101",--12169
"010010000111000000000000000000101111",--12170
"001011000000000001010000000100101111",--12171
"101001000000000001000000000000000011",--12172
"000101000000000000000010111111000101",--12173
"001011000000000001100000000100101111",--12174
"101001000000000001000000000000000010",--12175
"000101000000000000000010111111000101",--12176
"001011000000000001100000000100101111",--12177
"101001000000000001000000000000000001",--12178
"000101000000000000000010111111000101",--12179
"011111001111000000100000000000000111",--12180
"001111001100000000110000000000000000",--12181
"011010000111000000000000000000100011",--12182
"001111001010000001000000000000000011",--12183
"111110000110001001000001100000000000",--12184
"001011000000000000110000000100101111",--12185
"101001000000000001000000000000000001",--12186
"000101000000000000000010111111000101",--12187
"001111001100000001100000000000000000",--12188
"010010001101000000000000000000011100",--12189
"001111001100000001110000000000000001",--12190
"111110001110001000110001100000000000",--12191
"001111001100000001110000000000000010",--12192
"111110001110001001000010000000000000",--12193
"111110000110000001000001100000000000",--12194
"001111001100000001000000000000000011",--12195
"111110001000001001010010000000000000",--12196
"111110000110000001000001100000000000",--12197
"001111001010000001000000000000000011",--12198
"111110000110001000110010100000000000",--12199
"111110001100001001000010000000000000",--12200
"111110001010010001000010000000000000",--12201
"010110001001000000000000000000001111",--12202
"001101001000000001000000000000000110",--12203
"011100001001000000000000000000000110",--12204
"111110001000100000000010000000000000",--12205
"111110000110010001000001100000000000",--12206
"001111001100000001000000000000000100",--12207
"111110000110001001000001100000000000",--12208
"001011000000000000110000000100101111",--12209
"000101000000000000000010111110111000",--12210
"111110001000100000000010000000000000",--12211
"111110000110000001000001100000000000",--12212
"001111001100000001000000000000000100",--12213
"111110000110001001000001100000000000",--12214
"001011000000000000110000000100101111",--12215
"101001000000000001000000000000000001",--12216
"000101000000000000000010111111000101",--12217
"001101000110000000110000000101101101",--12218
"001101000110000000110000000000000110",--12219
"010000000111000000000000000001000010",--12220
"001101111100000000110000000000000000",--12221
"101001000000000000010000000000000001",--12222
"001001111100000111111111111111111011",--12223
"101001111100010111100000000000000110",--12224
"000111000000000000000010011110011001",--12225
"101001111100000111100000000000000110",--12226
"001101111100000111111111111111111011",--12227
"000101000000000000000010111111111111",--12228
"001111000000000000110000000100101111",--12229
"001001111100000000101111111111111011",--12230
"010110000111000000000000000000101111",--12231
"001111000000000001000000000100101101",--12232
"010110001001000000110000000000101101",--12233
"001101111100000001010000000000000000",--12234
"001101001010000001100000000000000000",--12235
"101111001001110001000011110000100011",--12236
"101111001001100001001101011100001010",--12237
"111110000110000001000001100000000000",--12238
"001111001100000001000000000000000000",--12239
"111110001000001000110010000000000000",--12240
"001111000000000001010000000100010010",--12241
"111110001000000001010010000000000000",--12242
"001111001100000001010000000000000001",--12243
"111110001010001000110010100000000000",--12244
"001111000000000001100000000100010011",--12245
"111110001010000001100010100000000000",--12246
"001111001100000001100000000000000010",--12247
"111110001100001000110011000000000000",--12248
"001111000000000001110000000100010100",--12249
"111110001100000001110011000000000000",--12250
"001001111100000001001111111111111010",--12251
"001001111100000000111111111111111001",--12252
"001011111100000001101111111111111000",--12253
"001011111100000001011111111111110111",--12254
"001011111100000001001111111111110110",--12255
"001011111100000000111111111111110101",--12256
"101000000001111000000000100000000000",--12257
"101110001001111000000001100000000000",--12258
"101110001011111000000010000000000000",--12259
"101110001101111000000010100000000000",--12260
"001001111100000111111111111111110100",--12261
"101001111100010111100000000000001101",--12262
"000111000000000000000000011110001000",--12263
"101001111100000111100000000000001101",--12264
"001101111100000111111111111111110100",--12265
"010000000011000000000000000000001100",--12266
"001111111100000000111111111111110101",--12267
"001011000000000000110000000100101101",--12268
"001111111100000000111111111111110110",--12269
"001011000000000000110000000100101010",--12270
"001111111100000000111111111111110111",--12271
"001011000000000000110000000100101011",--12272
"001111111100000000111111111111111000",--12273
"001011000000000000110000000100101100",--12274
"001101111100000000011111111111111001",--12275
"001001000000000000010000000100101001",--12276
"001101111100000000011111111111111010",--12277
"001001000000000000010000000100101110",--12278
"101001000000000000010000000000000001",--12279
"001101111100000000101111111111111011",--12280
"001101111100000000110000000000000000",--12281
"001001111100000111111111111111111010",--12282
"101001111100010111100000000000000111",--12283
"000111000000000000000010011110011001",--12284
"101001111100000111100000000000000111",--12285
"001101111100000111111111111111111010",--12286
"001101111100000000011111111111111100",--12287
"001101000010000000100000000000000011",--12288
"010011000101000000000000000000001110",--12289
"001101000100000000100000000100110001",--12290
"001101111100000000110000000000000000",--12291
"101000000001111000000000100000000000",--12292
"001001111100000111111111111111111011",--12293
"101001111100010111100000000000000110",--12294
"000111000000000000000010011110011001",--12295
"101001111100000111100000000000000110",--12296
"101001000000000000010000000000000100",--12297
"001101111100000000101111111111111100",--12298
"001101111100000000110000000000000000",--12299
"101001111100010111100000000000000110",--12300
"000111000000000000000010101111001101",--12301
"101001111100000111100000000000000110",--12302
"001101111100000111111111111111111011",--12303
"001101111100000000011111111111111110",--12304
"101001000010000000010000000000000001",--12305
"001101111100000000111111111111111111",--12306
"001100000110000000010001000000000000",--12307
"001101000100000001000000000000000000",--12308
"010011001000000000001111100000000000",--12309
"001001111100000000011111111111111101",--12310
"011111001001011000110000000011001001",--12311
"001101000100000001000000000000000001",--12312
"010011001001000000000000000111110101",--12313
"001101001000000001000000000100110001",--12314
"001101001000000001010000000000000000",--12315
"001001111100000000101111111111111100",--12316
"010011001011000000000000000010110001",--12317
"001101001010000001100000000101101101",--12318
"001101001100000001110000000000001010",--12319
"001111001110000000110000000000000000",--12320
"001111001110000001000000000000000001",--12321
"001111001110000001010000000000000010",--12322
"001101111100000010000000000000000000",--12323
"001101010000000010010000000000000001",--12324
"001100010010000001010100100000000000",--12325
"001101001100000010100000000000000001",--12326
"011111010101000000010000000000111011",--12327
"001101010000000001110000000000000000",--12328
"001111010010000001100000000000000000",--12329
"111110001100010000110011000000000000",--12330
"001111010010000001110000000000000001",--12331
"111110001100001001110011000000000000",--12332
"001111001110000001110000000000000001",--12333
"111110001100001001110011100000000000",--12334
"111110001110000001000011100000000001",--12335
"001101001100000001100000000000000100",--12336
"001111001100000010000000000000000001",--12337
"010110010001000001110000000000000111",--12338
"001111001110000001110000000000000010",--12339
"111110001100001001110011100000000000",--12340
"111110001110000001010011100000000001",--12341
"001111001100000010000000000000000010",--12342
"010110010001000001110000000000000010",--12343
"001111010010000001110000000000000001",--12344
"011110001111000000000000000000100110",--12345
"001111010010000001100000000000000010",--12346
"111110001100010001000011000000000000",--12347
"001111010010000001110000000000000011",--12348
"111110001100001001110011000000000000",--12349
"001111001110000001110000000000000000",--12350
"111110001100001001110011100000000000",--12351
"111110001110000000110011100000000001",--12352
"001111001100000010000000000000000000",--12353
"010110010001000001110000000000000111",--12354
"001111001110000001110000000000000010",--12355
"111110001100001001110011100000000000",--12356
"111110001110000001010011100000000001",--12357
"001111001100000010000000000000000010",--12358
"010110010001000001110000000000000010",--12359
"001111010010000001110000000000000011",--12360
"011110001111000000000000000000010011",--12361
"001111010010000001100000000000000100",--12362
"111110001100010001010010100000000000",--12363
"001111010010000001100000000000000101",--12364
"111110001010001001100010100000000000",--12365
"001111001110000001100000000000000000",--12366
"111110001010001001100011000000000000",--12367
"111110001100000000110001100000000001",--12368
"001111001100000001100000000000000000",--12369
"010110001101000000110000000000110110",--12370
"001111001110000000110000000000000001",--12371
"111110001010001000110001100000000000",--12372
"111110000110000001000001100000000001",--12373
"001111001100000001000000000000000001",--12374
"010110001001000000110000000000110001",--12375
"001111010010000000110000000000000101",--12376
"010010000111000000000000000000101111",--12377
"001011000000000001010000000100101111",--12378
"101001000000000001100000000000000011",--12379
"000101000000000000000011000010010101",--12380
"001011000000000001100000000100101111",--12381
"101001000000000001100000000000000010",--12382
"000101000000000000000011000010010101",--12383
"001011000000000001100000000100101111",--12384
"101001000000000001100000000000000001",--12385
"000101000000000000000011000010010101",--12386
"011111010101000000100000000000000111",--12387
"001111010010000000110000000000000000",--12388
"011010000111000000000000000000100011",--12389
"001111001110000001000000000000000011",--12390
"111110000110001001000001100000000000",--12391
"001011000000000000110000000100101111",--12392
"101001000000000001100000000000000001",--12393
"000101000000000000000011000010010101",--12394
"001111010010000001100000000000000000",--12395
"010010001101000000000000000000011100",--12396
"001111010010000001110000000000000001",--12397
"111110001110001000110001100000000000",--12398
"001111010010000001110000000000000010",--12399
"111110001110001001000010000000000000",--12400
"111110000110000001000001100000000000",--12401
"001111010010000001000000000000000011",--12402
"111110001000001001010010000000000000",--12403
"111110000110000001000001100000000000",--12404
"001111001110000001000000000000000011",--12405
"111110000110001000110010100000000000",--12406
"111110001100001001000010000000000000",--12407
"111110001010010001000010000000000000",--12408
"010110001001000000000000000000001111",--12409
"001101001100000001100000000000000110",--12410
"011100001101000000000000000000000110",--12411
"111110001000100000000010000000000000",--12412
"111110000110010001000001100000000000",--12413
"001111010010000001000000000000000100",--12414
"111110000110001001000001100000000000",--12415
"001011000000000000110000000100101111",--12416
"000101000000000000000011000010000111",--12417
"111110001000100000000010000000000000",--12418
"111110000110000001000001100000000000",--12419
"001111010010000001000000000000000100",--12420
"111110000110001001000001100000000000",--12421
"001011000000000000110000000100101111",--12422
"101001000000000001100000000000000001",--12423
"000101000000000000000011000010010101",--12424
"001101001010000001010000000101101101",--12425
"001101001010000001010000000000000110",--12426
"010000001011000000000000000001000011",--12427
"101000010001111000000001100000000000",--12428
"101000001001111000000001000000000000",--12429
"101001000000000000010000000000000001",--12430
"001001111100000111111111111111111011",--12431
"101001111100010111100000000000000110",--12432
"000111000000000000000010011110011001",--12433
"101001111100000111100000000000000110",--12434
"001101111100000111111111111111111011",--12435
"000101000000000000000011000011001111",--12436
"001111000000000000110000000100101111",--12437
"001001111100000001001111111111111011",--12438
"010110000111000000000000000000101111",--12439
"001111000000000001000000000100101101",--12440
"010110001001000000110000000000101101",--12441
"001101010000000001110000000000000000",--12442
"101111001001110001000011110000100011",--12443
"101111001001100001001101011100001010",--12444
"111110000110000001000001100000000000",--12445
"001111001110000001000000000000000000",--12446
"111110001000001000110010000000000000",--12447
"001111000000000001010000000100010010",--12448
"111110001000000001010010000000000000",--12449
"001111001110000001010000000000000001",--12450
"111110001010001000110010100000000000",--12451
"001111000000000001100000000100010011",--12452
"111110001010000001100010100000000000",--12453
"001111001110000001100000000000000010",--12454
"111110001100001000110011000000000000",--12455
"001111000000000001110000000100010100",--12456
"111110001100000001110011000000000000",--12457
"001001111100000001101111111111111010",--12458
"001001111100000001011111111111111001",--12459
"001011111100000001101111111111111000",--12460
"001011111100000001011111111111110111",--12461
"001011111100000001001111111111110110",--12462
"001011111100000000111111111111110101",--12463
"101000001001111000000001000000000000",--12464
"101000000001111000000000100000000000",--12465
"101110001001111000000001100000000000",--12466
"101110001011111000000010000000000000",--12467
"101110001101111000000010100000000000",--12468
"001001111100000111111111111111110100",--12469
"101001111100010111100000000000001101",--12470
"000111000000000000000000011110001000",--12471
"101001111100000111100000000000001101",--12472
"001101111100000111111111111111110100",--12473
"010000000011000000000000000000001100",--12474
"001111111100000000111111111111110101",--12475
"001011000000000000110000000100101101",--12476
"001111111100000000111111111111110110",--12477
"001011000000000000110000000100101010",--12478
"001111111100000000111111111111110111",--12479
"001011000000000000110000000100101011",--12480
"001111111100000000111111111111111000",--12481
"001011000000000000110000000100101100",--12482
"001101111100000000011111111111111001",--12483
"001001000000000000010000000100101001",--12484
"001101111100000000011111111111111010",--12485
"001001000000000000010000000100101110",--12486
"101001000000000000010000000000000001",--12487
"001101111100000000101111111111111011",--12488
"001101111100000000110000000000000000",--12489
"001001111100000111111111111111111010",--12490
"101001111100010111100000000000000111",--12491
"000111000000000000000010011110011001",--12492
"101001111100000111100000000000000111",--12493
"001101111100000111111111111111111010",--12494
"001101111100000000011111111111111100",--12495
"001101000010000000100000000000000010",--12496
"010011000101000000000000000100111101",--12497
"001101000100000000100000000100110001",--12498
"001101111100000000110000000000000000",--12499
"101000000001111000000000100000000000",--12500
"001001111100000111111111111111111011",--12501
"101001111100010111100000000000000110",--12502
"000111000000000000000010011110011001",--12503
"101001111100000111100000000000000110",--12504
"101001000000000000010000000000000011",--12505
"001101111100000000101111111111111100",--12506
"001101111100000000110000000000000000",--12507
"101001111100010111100000000000000110",--12508
"000111000000000000000010101111001101",--12509
"101001111100000111100000000000000110",--12510
"001101111100000111111111111111111011",--12511
"000101000000000000000011001000001111",--12512
"001101001000000001010000000101101101",--12513
"001101001010000001100000000000001010",--12514
"001111001100000000110000000000000000",--12515
"001111001100000001000000000000000001",--12516
"001111001100000001010000000000000010",--12517
"001101111100000001110000000000000000",--12518
"001101001110000010000000000000000001",--12519
"001100010000000001000010000000000000",--12520
"001101001010000010010000000000000001",--12521
"011111010011000000010000000000111000",--12522
"001101001110000001100000000000000000",--12523
"001111001000000001100000000000000000",--12524
"111110001100010000110011000000000000",--12525
"001111001000000001110000000000000001",--12526
"111110001100001001110011000000000000",--12527
"001111001100000001110000000000000001",--12528
"111110001100001001110011100000000000",--12529
"111110001110000001000011100000000001",--12530
"001101001010000001010000000000000100",--12531
"001111001010000010000000000000000001",--12532
"010110010001000001110000000000000111",--12533
"001111001100000001110000000000000010",--12534
"111110001100001001110011100000000000",--12535
"111110001110000001010011100000000001",--12536
"001111001010000010000000000000000010",--12537
"010110010001000001110000000000000010",--12538
"001111001000000001110000000000000001",--12539
"011110001111000000000000000000100100",--12540
"001111001000000001100000000000000010",--12541
"111110001100010001000011000000000000",--12542
"001111001000000001110000000000000011",--12543
"111110001100001001110011000000000000",--12544
"001111001100000001110000000000000000",--12545
"111110001100001001110011100000000000",--12546
"111110001110000000110011100000000001",--12547
"001111001010000010000000000000000000",--12548
"010110010001000001110000000000000111",--12549
"001111001100000001110000000000000010",--12550
"111110001100001001110011100000000000",--12551
"111110001110000001010011100000000001",--12552
"001111001010000010000000000000000010",--12553
"010110010001000001110000000000000010",--12554
"001111001000000001110000000000000011",--12555
"011110001111000000000000000000010010",--12556
"001111001000000001100000000000000100",--12557
"111110001100010001010010100000000000",--12558
"001111001000000001100000000000000101",--12559
"111110001010001001100010100000000000",--12560
"001111001100000001100000000000000000",--12561
"111110001010001001100011000000000000",--12562
"111110001100000000110001100000000001",--12563
"001111001010000001100000000000000000",--12564
"010110001101000000110000000011111001",--12565
"001111001100000000110000000000000001",--12566
"111110001010001000110001100000000000",--12567
"111110000110000001000001100000000001",--12568
"001111001010000001000000000000000001",--12569
"010110001001000000110000000011110100",--12570
"001111001000000000110000000000000101",--12571
"010010000111000000000000000011110010",--12572
"001011000000000001010000000100101111",--12573
"000101000000000000000011000101000110",--12574
"001011000000000001100000000100101111",--12575
"000101000000000000000011000101000110",--12576
"001011000000000001100000000100101111",--12577
"000101000000000000000011000101000110",--12578
"011111010011000000100000000000000110",--12579
"001111001000000000110000000000000000",--12580
"011010000111000000000000000011101001",--12581
"001111001100000001000000000000000011",--12582
"111110000110001001000001100000000000",--12583
"001011000000000000110000000100101111",--12584
"000101000000000000000011000101000110",--12585
"001111001000000001100000000000000000",--12586
"010010001101000000000000000011100011",--12587
"001111001000000001110000000000000001",--12588
"111110001110001000110001100000000000",--12589
"001111001000000001110000000000000010",--12590
"111110001110001001000010000000000000",--12591
"111110000110000001000001100000000000",--12592
"001111001000000001000000000000000011",--12593
"111110001000001001010010000000000000",--12594
"111110000110000001000001100000000000",--12595
"001111001100000001000000000000000011",--12596
"111110000110001000110010100000000000",--12597
"111110001100001001000010000000000000",--12598
"111110001010010001000010000000000000",--12599
"010110001001000000000000000011010110",--12600
"001101001010000001010000000000000110",--12601
"011100001011000000000000000000000110",--12602
"111110001000100000000010000000000000",--12603
"111110000110010001000001100000000000",--12604
"001111001000000001000000000000000100",--12605
"111110000110001001000001100000000000",--12606
"001011000000000000110000000100101111",--12607
"000101000000000000000011000101000110",--12608
"111110001000100000000010000000000000",--12609
"111110000110000001000001100000000000",--12610
"001111001000000001000000000000000100",--12611
"111110000110001001000001100000000000",--12612
"001011000000000000110000000100101111",--12613
"001111000000000000110000000100101111",--12614
"001111000000000001000000000100101101",--12615
"010110001001000000110000000011000110",--12616
"001101000100000001000000000000000001",--12617
"010011001001000000000000000011000100",--12618
"001101001000000001000000000100110001",--12619
"001101001000000001010000000000000000",--12620
"001001111100000000101111111111111100",--12621
"010011001011000000000000000010101111",--12622
"001101001010000001100000000101101101",--12623
"001101001100000010010000000000001010",--12624
"001111010010000000110000000000000000",--12625
"001111010010000001000000000000000001",--12626
"001111010010000001010000000000000010",--12627
"001100010000000001010100000000000000",--12628
"001101001100000010100000000000000001",--12629
"011111010101000000010000000000111011",--12630
"001101001110000010010000000000000000",--12631
"001111010000000001100000000000000000",--12632
"111110001100010000110011000000000000",--12633
"001111010000000001110000000000000001",--12634
"111110001100001001110011000000000000",--12635
"001111010010000001110000000000000001",--12636
"111110001100001001110011100000000000",--12637
"111110001110000001000011100000000001",--12638
"001101001100000001100000000000000100",--12639
"001111001100000010000000000000000001",--12640
"010110010001000001110000000000000111",--12641
"001111010010000001110000000000000010",--12642
"111110001100001001110011100000000000",--12643
"111110001110000001010011100000000001",--12644
"001111001100000010000000000000000010",--12645
"010110010001000001110000000000000010",--12646
"001111010000000001110000000000000001",--12647
"011110001111000000000000000000100110",--12648
"001111010000000001100000000000000010",--12649
"111110001100010001000011000000000000",--12650
"001111010000000001110000000000000011",--12651
"111110001100001001110011000000000000",--12652
"001111010010000001110000000000000000",--12653
"111110001100001001110011100000000000",--12654
"111110001110000000110011100000000001",--12655
"001111001100000010000000000000000000",--12656
"010110010001000001110000000000000111",--12657
"001111010010000001110000000000000010",--12658
"111110001100001001110011100000000000",--12659
"111110001110000001010011100000000001",--12660
"001111001100000010000000000000000010",--12661
"010110010001000001110000000000000010",--12662
"001111010000000001110000000000000011",--12663
"011110001111000000000000000000010011",--12664
"001111010000000001100000000000000100",--12665
"111110001100010001010010100000000000",--12666
"001111010000000001100000000000000101",--12667
"111110001010001001100010100000000000",--12668
"001111010010000001100000000000000000",--12669
"111110001010001001100011000000000000",--12670
"111110001100000000110001100000000001",--12671
"001111001100000001100000000000000000",--12672
"010110001101000000110000000000110110",--12673
"001111010010000000110000000000000001",--12674
"111110001010001000110001100000000000",--12675
"111110000110000001000001100000000001",--12676
"001111001100000001000000000000000001",--12677
"010110001001000000110000000000110001",--12678
"001111010000000000110000000000000101",--12679
"010010000111000000000000000000101111",--12680
"001011000000000001010000000100101111",--12681
"101001000000000001100000000000000011",--12682
"000101000000000000000011000111000100",--12683
"001011000000000001100000000100101111",--12684
"101001000000000001100000000000000010",--12685
"000101000000000000000011000111000100",--12686
"001011000000000001100000000100101111",--12687
"101001000000000001100000000000000001",--12688
"000101000000000000000011000111000100",--12689
"011111010101000000100000000000000111",--12690
"001111010000000000110000000000000000",--12691
"011010000111000000000000000000100011",--12692
"001111010010000001000000000000000011",--12693
"111110000110001001000001100000000000",--12694
"001011000000000000110000000100101111",--12695
"101001000000000001100000000000000001",--12696
"000101000000000000000011000111000100",--12697
"001111010000000001100000000000000000",--12698
"010010001101000000000000000000011100",--12699
"001111010000000001110000000000000001",--12700
"111110001110001000110001100000000000",--12701
"001111010000000001110000000000000010",--12702
"111110001110001001000010000000000000",--12703
"111110000110000001000001100000000000",--12704
"001111010000000001000000000000000011",--12705
"111110001000001001010010000000000000",--12706
"111110000110000001000001100000000000",--12707
"001111010010000001000000000000000011",--12708
"111110000110001000110010100000000000",--12709
"111110001100001001000010000000000000",--12710
"111110001010010001000010000000000000",--12711
"010110001001000000000000000000001111",--12712
"001101001100000001100000000000000110",--12713
"011100001101000000000000000000000110",--12714
"111110001000100000000010000000000000",--12715
"111110000110010001000001100000000000",--12716
"001111010000000001000000000000000100",--12717
"111110000110001001000001100000000000",--12718
"001011000000000000110000000100101111",--12719
"000101000000000000000011000110110110",--12720
"111110001000100000000010000000000000",--12721
"111110000110000001000001100000000000",--12722
"001111010000000001000000000000000100",--12723
"111110000110001001000001100000000000",--12724
"001011000000000000110000000100101111",--12725
"101001000000000001100000000000000001",--12726
"000101000000000000000011000111000100",--12727
"001101001010000001010000000101101101",--12728
"001101001010000001010000000000000110",--12729
"010000001011000000000000000001000011",--12730
"101000001111111000000001100000000000",--12731
"101000001001111000000001000000000000",--12732
"101001000000000000010000000000000001",--12733
"001001111100000111111111111111111011",--12734
"101001111100010111100000000000000110",--12735
"000111000000000000000010011110011001",--12736
"101001111100000111100000000000000110",--12737
"001101111100000111111111111111111011",--12738
"000101000000000000000011000111111110",--12739
"001111000000000000110000000100101111",--12740
"001001111100000001001111111111111011",--12741
"010110000111000000000000000000101111",--12742
"001111000000000001000000000100101101",--12743
"010110001001000000110000000000101101",--12744
"001101001110000010000000000000000000",--12745
"101111001001110001000011110000100011",--12746
"101111001001100001001101011100001010",--12747
"111110000110000001000001100000000000",--12748
"001111010000000001000000000000000000",--12749
"111110001000001000110010000000000000",--12750
"001111000000000001010000000100010010",--12751
"111110001000000001010010000000000000",--12752
"001111010000000001010000000000000001",--12753
"111110001010001000110010100000000000",--12754
"001111000000000001100000000100010011",--12755
"111110001010000001100010100000000000",--12756
"001111010000000001100000000000000010",--12757
"111110001100001000110011000000000000",--12758
"001111000000000001110000000100010100",--12759
"111110001100000001110011000000000000",--12760
"001001111100000001101111111111111010",--12761
"001001111100000001011111111111111001",--12762
"001011111100000001101111111111111000",--12763
"001011111100000001011111111111110111",--12764
"001011111100000001001111111111110110",--12765
"001011111100000000111111111111110101",--12766
"101000001001111000000001000000000000",--12767
"101000000001111000000000100000000000",--12768
"101110001001111000000001100000000000",--12769
"101110001011111000000010000000000000",--12770
"101110001101111000000010100000000000",--12771
"001001111100000111111111111111110100",--12772
"101001111100010111100000000000001101",--12773
"000111000000000000000000011110001000",--12774
"101001111100000111100000000000001101",--12775
"001101111100000111111111111111110100",--12776
"010000000011000000000000000000001100",--12777
"001111111100000000111111111111110101",--12778
"001011000000000000110000000100101101",--12779
"001111111100000000111111111111110110",--12780
"001011000000000000110000000100101010",--12781
"001111111100000000111111111111110111",--12782
"001011000000000000110000000100101011",--12783
"001111111100000000111111111111111000",--12784
"001011000000000000110000000100101100",--12785
"001101111100000000011111111111111001",--12786
"001001000000000000010000000100101001",--12787
"001101111100000000011111111111111010",--12788
"001001000000000000010000000100101110",--12789
"101001000000000000010000000000000001",--12790
"001101111100000000101111111111111011",--12791
"001101111100000000110000000000000000",--12792
"001001111100000111111111111111111010",--12793
"101001111100010111100000000000000111",--12794
"000111000000000000000010011110011001",--12795
"101001111100000111100000000000000111",--12796
"001101111100000111111111111111111010",--12797
"001101111100000000011111111111111100",--12798
"001101000010000000100000000000000010",--12799
"010011000101000000000000000000001110",--12800
"001101000100000000100000000100110001",--12801
"001101111100000000110000000000000000",--12802
"101000000001111000000000100000000000",--12803
"001001111100000111111111111111111011",--12804
"101001111100010111100000000000000110",--12805
"000111000000000000000010011110011001",--12806
"101001111100000111100000000000000110",--12807
"101001000000000000010000000000000011",--12808
"001101111100000000101111111111111100",--12809
"001101111100000000110000000000000000",--12810
"101001111100010111100000000000000110",--12811
"000111000000000000000010101111001101",--12812
"101001111100000111100000000000000110",--12813
"001101111100000111111111111111111011",--12814
"001101111100000000011111111111111101",--12815
"101001000010000000010000000000000001",--12816
"001101111100000000101111111111111111",--12817
"001101111100000000110000000000000000",--12818
"000101000000000000000010110111111111",--12819
"010111000010000000001111100000000000",--12820
"001101000010000000110000000000000100",--12821
"001101000110000001000000000000000001",--12822
"101111001011110001010100111001101110",--12823
"101111001011100001010110101100101000",--12824
"001011000000000001010000000100101101",--12825
"001101000000000001100000000100110000",--12826
"001001111100000000010000000000000000",--12827
"001011111100000001001111111111111111",--12828
"001001111100000000101111111111111110",--12829
"001011111100000000111111111111111101",--12830
"001001111100000001001111111111111100",--12831
"001001111100000000111111111111111011",--12832
"101000001001111000000001100000000000",--12833
"101000001101111000000001000000000000",--12834
"101000000001111000000000100000000000",--12835
"001001111100000111111111111111111010",--12836
"101001111100010111100000000000000111",--12837
"000111000000000000000010110111111111",--12838
"101001111100000111100000000000000111",--12839
"001101111100000111111111111111111010",--12840
"001111000000000000110000000100101101",--12841
"101111001001110001001011110111001100",--12842
"101111001001100001001100110011001101",--12843
"010110000111000001000000001010111001",--12844
"101111001001110001000100110010111110",--12845
"101111001001100001001011110000100000",--12846
"010110001001000000110000001010110110",--12847
"001101000000000000010000000100101001",--12848
"101000000011000000010000100010000010",--12849
"001101000000000000100000000100101110",--12850
"101000000010000000100000100000000000",--12851
"001101111100000000101111111111111011",--12852
"001101000100000000110000000000000000",--12853
"011100000011000000110000001010101111",--12854
"001101000000000000010000000100110000",--12855
"001101000010000000110000000000000000",--12856
"001101000110000001000000000000000000",--12857
"010011001001000000000000001001101110",--12858
"001001111100000000111111111111111010",--12859
"001001111100000000011111111111111001",--12860
"010011001001011000110000000101111111",--12861
"001101001000000001010000000101101101",--12862
"001111000000000000110000000100101010",--12863
"001101001010000001100000000000000101",--12864
"001111001100000001000000000000000000",--12865
"111110000110010001000001100000000000",--12866
"001111000000000001000000000100101011",--12867
"001111001100000001010000000000000001",--12868
"111110001000010001010010000000000000",--12869
"001111000000000001010000000100101100",--12870
"001111001100000001100000000000000010",--12871
"111110001010010001100010100000000000",--12872
"001101001000000001000000000010111110",--12873
"001101001010000001100000000000000001",--12874
"011111001101000000010000000000110111",--12875
"001111001000000001100000000000000000",--12876
"111110001100010000110011000000000000",--12877
"001111001000000001110000000000000001",--12878
"111110001100001001110011000000000000",--12879
"001111000000000001110000000011111011",--12880
"111110001100001001110011100000000000",--12881
"111110001110000001000011100000000001",--12882
"001101001010000001010000000000000100",--12883
"001111001010000010000000000000000001",--12884
"010110010001000001110000000000000111",--12885
"001111000000000001110000000011111100",--12886
"111110001100001001110011100000000000",--12887
"111110001110000001010011100000000001",--12888
"001111001010000010000000000000000010",--12889
"010110010001000001110000000000000010",--12890
"001111001000000001110000000000000001",--12891
"011110001111000000000000000000100100",--12892
"001111001000000001100000000000000010",--12893
"111110001100010001000011000000000000",--12894
"001111001000000001110000000000000011",--12895
"111110001100001001110011000000000000",--12896
"001111000000000001110000000011111010",--12897
"111110001100001001110011100000000000",--12898
"111110001110000000110011100000000001",--12899
"001111001010000010000000000000000000",--12900
"010110010001000001110000000000000111",--12901
"001111000000000001110000000011111100",--12902
"111110001100001001110011100000000000",--12903
"111110001110000001010011100000000001",--12904
"001111001010000010000000000000000010",--12905
"010110010001000001110000000000000010",--12906
"001111001000000001110000000000000011",--12907
"011110001111000000000000000000010010",--12908
"001111001000000001100000000000000100",--12909
"111110001100010001010010100000000000",--12910
"001111001000000001100000000000000101",--12911
"111110001010001001100010100000000000",--12912
"001111000000000001100000000011111010",--12913
"111110001010001001100011000000000000",--12914
"111110001100000000110001100000000001",--12915
"001111001010000001100000000000000000",--12916
"010110001101000000110000000100111110",--12917
"001111000000000000110000000011111011",--12918
"111110001010001000110001100000000000",--12919
"111110000110000001000001100000000001",--12920
"001111001010000001000000000000000001",--12921
"010110001001000000110000000100111001",--12922
"001111001000000000110000000000000101",--12923
"010010000111000000000000000100110111",--12924
"001011000000000001010000000100101111",--12925
"000101000000000000000011001011001011",--12926
"001011000000000001100000000100101111",--12927
"000101000000000000000011001011001011",--12928
"001011000000000001100000000100101111",--12929
"000101000000000000000011001011001011",--12930
"011111001101000000100000000000001100",--12931
"001111001000000001100000000000000000",--12932
"011010001101000000000000000100101110",--12933
"001111001000000001100000000000000001",--12934
"111110001100001000110001100000000000",--12935
"001111001000000001100000000000000010",--12936
"111110001100001001000010000000000000",--12937
"111110000110000001000001100000000000",--12938
"001111001000000001000000000000000011",--12939
"111110001000001001010010000000000000",--12940
"111110000110000001000001100000000000",--12941
"001011000000000000110000000100101111",--12942
"000101000000000000000011001011001011",--12943
"001111001000000001100000000000000000",--12944
"010010001101000000000000000100100010",--12945
"001111001000000001110000000000000001",--12946
"111110001110001000110011100000000000",--12947
"001111001000000010000000000000000010",--12948
"111110010000001001000100000000000000",--12949
"111110001110000010000011100000000000",--12950
"001111001000000010000000000000000011",--12951
"111110010000001001010100000000000000",--12952
"111110001110000010000011100000000000",--12953
"111110000110001000110100000000000000",--12954
"001101001010000001110000000000000100",--12955
"001111001110000010010000000000000000",--12956
"111110010000001010010100000000000000",--12957
"111110001000001001000100100000000000",--12958
"001111001110000010100000000000000001",--12959
"111110010010001010100100100000000000",--12960
"111110010000000010010100000000000000",--12961
"111110001010001001010100100000000000",--12962
"001111001110000010100000000000000010",--12963
"111110010010001010100100100000000000",--12964
"111110010000000010010100000000000000",--12965
"001101001010000001110000000000000011",--12966
"011100001111000000000000000000000011",--12967
"101110010001111000000001100000000000",--12968
"011111001101000000110000000000010000",--12969
"000101000000000000000011001010111001",--12970
"111110001000001001010100100000000000",--12971
"001101001010000001110000000000001001",--12972
"001111001110000010100000000000000000",--12973
"111110010010001010100100100000000000",--12974
"111110010000000010010100000000000000",--12975
"111110001010001000110010100000000000",--12976
"001111001110000010010000000000000001",--12977
"111110001010001010010010100000000000",--12978
"111110010000000001010010100000000000",--12979
"111110000110001001000001100000000000",--12980
"001111001110000001000000000000000010",--12981
"111110000110001001000001100000000000",--12982
"111110001010000000110001100000000000",--12983
"011111001101000000110000000000000001",--12984
"111110000110010000010001100000000000",--12985
"111110001110001001110010000000000000",--12986
"111110001100001000110001100000000000",--12987
"111110001000010000110001100000000000",--12988
"010110000111000000000000000011110110",--12989
"001101001010000001010000000000000110",--12990
"011100001011000000000000000000000110",--12991
"111110000110100000000001100000000000",--12992
"111110001110010000110001100000000000",--12993
"001111001000000001000000000000000100",--12994
"111110000110001001000001100000000000",--12995
"001011000000000000110000000100101111",--12996
"000101000000000000000011001011001011",--12997
"111110000110100000000001100000000000",--12998
"111110001110000000110001100000000000",--12999
"001111001000000001000000000000000100",--13000
"111110000110001001000001100000000000",--13001
"001011000000000000110000000100101111",--13002
"001111000000000000110000000100101111",--13003
"101111001001110001001011110111001100",--13004
"101111001001100001001100110011001101",--13005
"010110001001000000110000000011100101",--13006
"001101000110000001000000000000000001",--13007
"010011001001000000000000000011100011",--13008
"001101001000000001000000000100110001",--13009
"001101001000000001010000000000000000",--13010
"010011001011000000000000000011001110",--13011
"001101001010000001100000000101101101",--13012
"001111000000000000110000000100101010",--13013
"001101001100000001110000000000000101",--13014
"001111001110000001000000000000000000",--13015
"111110000110010001000001100000000000",--13016
"001111000000000001000000000100101011",--13017
"001111001110000001010000000000000001",--13018
"111110001000010001010010000000000000",--13019
"001111000000000001010000000100101100",--13020
"001111001110000001100000000000000010",--13021
"111110001010010001100010100000000000",--13022
"001101001010000001110000000010111110",--13023
"001101001100000010000000000000000001",--13024
"011111010001000000010000000000111100",--13025
"001111001110000001100000000000000000",--13026
"111110001100010000110011000000000000",--13027
"001111001110000001110000000000000001",--13028
"111110001100001001110011000000000000",--13029
"001111000000000001110000000011111011",--13030
"111110001100001001110011100000000000",--13031
"111110001110000001000011100000000001",--13032
"001101001100000001100000000000000100",--13033
"001111001100000010000000000000000001",--13034
"010110010001000001110000000000000111",--13035
"001111000000000001110000000011111100",--13036
"111110001100001001110011100000000000",--13037
"111110001110000001010011100000000001",--13038
"001111001100000010000000000000000010",--13039
"010110010001000001110000000000000010",--13040
"001111001110000001110000000000000001",--13041
"011110001111000000000000000000101000",--13042
"001111001110000001100000000000000010",--13043
"111110001100010001000011000000000000",--13044
"001111001110000001110000000000000011",--13045
"111110001100001001110011000000000000",--13046
"001111000000000001110000000011111010",--13047
"111110001100001001110011100000000000",--13048
"111110001110000000110011100000000001",--13049
"001111001100000010000000000000000000",--13050
"010110010001000001110000000000000111",--13051
"001111000000000001110000000011111100",--13052
"111110001100001001110011100000000000",--13053
"111110001110000001010011100000000001",--13054
"001111001100000010000000000000000010",--13055
"010110010001000001110000000000000010",--13056
"001111001110000001110000000000000011",--13057
"011110001111000000000000000000010101",--13058
"001111001110000001100000000000000100",--13059
"111110001100010001010010100000000000",--13060
"001111001110000001100000000000000101",--13061
"111110001010001001100010100000000000",--13062
"001111000000000001100000000011111010",--13063
"111110001010001001100011000000000000",--13064
"111110001100000000110001100000000001",--13065
"001111001100000001100000000000000000",--13066
"010110001101000000110000000000000111",--13067
"001111000000000000110000000011111011",--13068
"111110001010001000110001100000000000",--13069
"111110000110000001000001100000000001",--13070
"001111001100000001000000000000000001",--13071
"010110001001000000110000000000000010",--13072
"001111001110000000110000000000000101",--13073
"011110000111000000000000000000000010",--13074
"101000000001111000000011000000000000",--13075
"000101000000000000000011001101101110",--13076
"001011000000000001010000000100101111",--13077
"101001000000000001100000000000000011",--13078
"000101000000000000000011001101101110",--13079
"001011000000000001100000000100101111",--13080
"101001000000000001100000000000000010",--13081
"000101000000000000000011001101101110",--13082
"001011000000000001100000000100101111",--13083
"101001000000000001100000000000000001",--13084
"000101000000000000000011001101101110",--13085
"011111010001000000100000000000001111",--13086
"001111001110000001100000000000000000",--13087
"011010001101000000000000000000001011",--13088
"001111001110000001100000000000000001",--13089
"111110001100001000110001100000000000",--13090
"001111001110000001100000000000000010",--13091
"111110001100001001000010000000000000",--13092
"111110000110000001000001100000000000",--13093
"001111001110000001000000000000000011",--13094
"111110001000001001010010000000000000",--13095
"111110000110000001000001100000000000",--13096
"001011000000000000110000000100101111",--13097
"101001000000000001100000000000000001",--13098
"000101000000000000000011001101101110",--13099
"101000000001111000000011000000000000",--13100
"000101000000000000000011001101101110",--13101
"001111001110000001100000000000000000",--13102
"011110001101000000000000000000000010",--13103
"101000000001111000000011000000000000",--13104
"000101000000000000000011001101101110",--13105
"001111001110000001110000000000000001",--13106
"111110001110001000110011100000000000",--13107
"001111001110000010000000000000000010",--13108
"111110010000001001000100000000000000",--13109
"111110001110000010000011100000000000",--13110
"001111001110000010000000000000000011",--13111
"111110010000001001010100000000000000",--13112
"111110001110000010000011100000000000",--13113
"111110000110001000110100000000000000",--13114
"001101001100000010010000000000000100",--13115
"001111010010000010010000000000000000",--13116
"111110010000001010010100000000000000",--13117
"111110001000001001000100100000000000",--13118
"001111010010000010100000000000000001",--13119
"111110010010001010100100100000000000",--13120
"111110010000000010010100000000000000",--13121
"111110001010001001010100100000000000",--13122
"001111010010000010100000000000000010",--13123
"111110010010001010100100100000000000",--13124
"111110010000000010010100000000000000",--13125
"001101001100000010010000000000000011",--13126
"011100010011000000000000000000000011",--13127
"101110010001111000000001100000000000",--13128
"011111010001000000110000000000010000",--13129
"000101000000000000000011001101011001",--13130
"111110001000001001010100100000000000",--13131
"001101001100000010010000000000001001",--13132
"001111010010000010100000000000000000",--13133
"111110010010001010100100100000000000",--13134
"111110010000000010010100000000000000",--13135
"111110001010001000110010100000000000",--13136
"001111010010000010010000000000000001",--13137
"111110001010001010010010100000000000",--13138
"111110010000000001010010100000000000",--13139
"111110000110001001000001100000000000",--13140
"001111010010000001000000000000000010",--13141
"111110000110001001000001100000000000",--13142
"111110001010000000110001100000000000",--13143
"011111010001000000110000000000000001",--13144
"111110000110010000010001100000000000",--13145
"111110001110001001110010000000000000",--13146
"111110001100001000110001100000000000",--13147
"111110001000010000110001100000000000",--13148
"010110000111000000000000000000001111",--13149
"001101001100000001100000000000000110",--13150
"011100001101000000000000000000000110",--13151
"111110000110100000000001100000000000",--13152
"111110001110010000110001100000000000",--13153
"001111001110000001000000000000000100",--13154
"111110000110001001000001100000000000",--13155
"001011000000000000110000000100101111",--13156
"000101000000000000000011001101101011",--13157
"111110000110100000000001100000000000",--13158
"111110001110000000110001100000000000",--13159
"001111001110000001000000000000000100",--13160
"111110000110001001000001100000000000",--13161
"001011000000000000110000000100101111",--13162
"101001000000000001100000000000000001",--13163
"000101000000000000000011001101101110",--13164
"101000000001111000000011000000000000",--13165
"001111000000000000110000000100101111",--13166
"010000001101000000000000000000100111",--13167
"101111001001110001001011111001001100",--13168
"101111001001100001001100110011001101",--13169
"010110001001000000110000000000100100",--13170
"101111001001110001000011110000100011",--13171
"101111001001100001001101011100001010",--13172
"111110000110000001000001100000000000",--13173
"001111000000000001000000000101100100",--13174
"111110001000001000110010000000000000",--13175
"001111000000000001010000000100101010",--13176
"111110001000000001010010000000000000",--13177
"001111000000000001010000000101100101",--13178
"111110001010001000110010100000000000",--13179
"001111000000000001100000000100101011",--13180
"111110001010000001100010100000000000",--13181
"001111000000000001100000000101100110",--13182
"111110001100001000110001100000000000",--13183
"001111000000000001100000000100101100",--13184
"111110000110000001100001100000000000",--13185
"001001111100000001001111111111111000",--13186
"101000001001111000000001000000000000",--13187
"101000000001111000000000100000000000",--13188
"101110001011111000001111100000000000",--13189
"101110000111111000000010100000000000",--13190
"101110001001111000000001100000000000",--13191
"101110111111111000000010000000000000",--13192
"001001111100000111111111111111110111",--13193
"101001111100010111100000000000001010",--13194
"000111000000000000000000011110001000",--13195
"101001111100000111100000000000001010",--13196
"001101111100000111111111111111110111",--13197
"011100000011000000000000000000101110",--13198
"101001000000000000010000000000000001",--13199
"001101111100000000101111111111111000",--13200
"101001111100010111100000000000001010",--13201
"000111000000000000000000100011100001",--13202
"101001111100000111100000000000001010",--13203
"001101111100000111111111111111110111",--13204
"011100000011000000000000000000100111",--13205
"000101000000000000000011001110100010",--13206
"001101001010000001010000000101101101",--13207
"001101001010000001010000000000000110",--13208
"010000001011000000000000000000001000",--13209
"101000001001111000000001000000000000",--13210
"101001000000000000010000000000000001",--13211
"001001111100000111111111111111111000",--13212
"101001111100010111100000000000001001",--13213
"000111000000000000000000100011100001",--13214
"101001111100000111100000000000001001",--13215
"001101111100000111111111111111111000",--13216
"011100000011000000000000000000011011",--13217
"001101111100000000011111111111111010",--13218
"001101000010000000100000000000000010",--13219
"010011000101000000000000000000001111",--13220
"001101000100000000100000000100110001",--13221
"101000000001111000000000100000000000",--13222
"001001111100000111111111111111111000",--13223
"101001111100010111100000000000001001",--13224
"000111000000000000000000100011100001",--13225
"101001111100000111100000000000001001",--13226
"001101111100000111111111111111111000",--13227
"011100000011000000000000000000010000",--13228
"101001000000000000010000000000000011",--13229
"001101111100000000101111111111111010",--13230
"101001111100010111100000000000001001",--13231
"000111000000000000000000110101111110",--13232
"101001111100000111100000000000001001",--13233
"001101111100000111111111111111111000",--13234
"011100000011000000000000000000001001",--13235
"101001000000000000010000000000000001",--13236
"001101111100000000101111111111111001",--13237
"001001111100000111111111111111111000",--13238
"101001111100010111100000000000001001",--13239
"000111000000000000000000111111111011",--13240
"101001111100000111100000000000001001",--13241
"001101111100000111111111111111111000",--13242
"011100000011000000000000000100101010",--13243
"000101000000000000000011010010101001",--13244
"001101111100000000011111111111111010",--13245
"001101000010000000100000000000000001",--13246
"010011000101000000000000000011100001",--13247
"001101000100000000100000000100110001",--13248
"001101000100000000110000000000000000",--13249
"010011000111000000000000000011001100",--13250
"001101000110000001000000000101101101",--13251
"001111000000000000110000000100101010",--13252
"001101001000000001010000000000000101",--13253
"001111001010000001000000000000000000",--13254
"111110000110010001000001100000000000",--13255
"001111000000000001000000000100101011",--13256
"001111001010000001010000000000000001",--13257
"111110001000010001010010000000000000",--13258
"001111000000000001010000000100101100",--13259
"001111001010000001100000000000000010",--13260
"111110001010010001100010100000000000",--13261
"001101000110000001010000000010111110",--13262
"001101001000000001100000000000000001",--13263
"011111001101000000010000000000111100",--13264
"001111001010000001100000000000000000",--13265
"111110001100010000110011000000000000",--13266
"001111001010000001110000000000000001",--13267
"111110001100001001110011000000000000",--13268
"001111000000000001110000000011111011",--13269
"111110001100001001110011100000000000",--13270
"111110001110000001000011100000000001",--13271
"001101001000000001000000000000000100",--13272
"001111001000000010000000000000000001",--13273
"010110010001000001110000000000000111",--13274
"001111000000000001110000000011111100",--13275
"111110001100001001110011100000000000",--13276
"111110001110000001010011100000000001",--13277
"001111001000000010000000000000000010",--13278
"010110010001000001110000000000000010",--13279
"001111001010000001110000000000000001",--13280
"011110001111000000000000000000101000",--13281
"001111001010000001100000000000000010",--13282
"111110001100010001000011000000000000",--13283
"001111001010000001110000000000000011",--13284
"111110001100001001110011000000000000",--13285
"001111000000000001110000000011111010",--13286
"111110001100001001110011100000000000",--13287
"111110001110000000110011100000000001",--13288
"001111001000000010000000000000000000",--13289
"010110010001000001110000000000000111",--13290
"001111000000000001110000000011111100",--13291
"111110001100001001110011100000000000",--13292
"111110001110000001010011100000000001",--13293
"001111001000000010000000000000000010",--13294
"010110010001000001110000000000000010",--13295
"001111001010000001110000000000000011",--13296
"011110001111000000000000000000010101",--13297
"001111001010000001100000000000000100",--13298
"111110001100010001010010100000000000",--13299
"001111001010000001100000000000000101",--13300
"111110001010001001100010100000000000",--13301
"001111000000000001100000000011111010",--13302
"111110001010001001100011000000000000",--13303
"111110001100000000110001100000000001",--13304
"001111001000000001100000000000000000",--13305
"010110001101000000110000000000000111",--13306
"001111000000000000110000000011111011",--13307
"111110001010001000110001100000000000",--13308
"111110000110000001000001100000000001",--13309
"001111001000000001000000000000000001",--13310
"010110001001000000110000000000000010",--13311
"001111001010000000110000000000000101",--13312
"011110000111000000000000000000000010",--13313
"101000000001111000000010000000000000",--13314
"000101000000000000000011010001011101",--13315
"001011000000000001010000000100101111",--13316
"101001000000000001000000000000000011",--13317
"000101000000000000000011010001011101",--13318
"001011000000000001100000000100101111",--13319
"101001000000000001000000000000000010",--13320
"000101000000000000000011010001011101",--13321
"001011000000000001100000000100101111",--13322
"101001000000000001000000000000000001",--13323
"000101000000000000000011010001011101",--13324
"011111001101000000100000000000001111",--13325
"001111001010000001100000000000000000",--13326
"011010001101000000000000000000001011",--13327
"001111001010000001100000000000000001",--13328
"111110001100001000110001100000000000",--13329
"001111001010000001100000000000000010",--13330
"111110001100001001000010000000000000",--13331
"111110000110000001000001100000000000",--13332
"001111001010000001000000000000000011",--13333
"111110001000001001010010000000000000",--13334
"111110000110000001000001100000000000",--13335
"001011000000000000110000000100101111",--13336
"101001000000000001000000000000000001",--13337
"000101000000000000000011010001011101",--13338
"101000000001111000000010000000000000",--13339
"000101000000000000000011010001011101",--13340
"001111001010000001100000000000000000",--13341
"011110001101000000000000000000000010",--13342
"101000000001111000000010000000000000",--13343
"000101000000000000000011010001011101",--13344
"001111001010000001110000000000000001",--13345
"111110001110001000110011100000000000",--13346
"001111001010000010000000000000000010",--13347
"111110010000001001000100000000000000",--13348
"111110001110000010000011100000000000",--13349
"001111001010000010000000000000000011",--13350
"111110010000001001010100000000000000",--13351
"111110001110000010000011100000000000",--13352
"111110000110001000110100000000000000",--13353
"001101001000000001110000000000000100",--13354
"001111001110000010010000000000000000",--13355
"111110010000001010010100000000000000",--13356
"111110001000001001000100100000000000",--13357
"001111001110000010100000000000000001",--13358
"111110010010001010100100100000000000",--13359
"111110010000000010010100000000000000",--13360
"111110001010001001010100100000000000",--13361
"001111001110000010100000000000000010",--13362
"111110010010001010100100100000000000",--13363
"111110010000000010010100000000000000",--13364
"001101001000000001110000000000000011",--13365
"011100001111000000000000000000000011",--13366
"101110010001111000000001100000000000",--13367
"011111001101000000110000000000010000",--13368
"000101000000000000000011010001001000",--13369
"111110001000001001010100100000000000",--13370
"001101001000000001110000000000001001",--13371
"001111001110000010100000000000000000",--13372
"111110010010001010100100100000000000",--13373
"111110010000000010010100000000000000",--13374
"111110001010001000110010100000000000",--13375
"001111001110000010010000000000000001",--13376
"111110001010001010010010100000000000",--13377
"111110010000000001010010100000000000",--13378
"111110000110001001000001100000000000",--13379
"001111001110000001000000000000000010",--13380
"111110000110001001000001100000000000",--13381
"111110001010000000110001100000000000",--13382
"011111001101000000110000000000000001",--13383
"111110000110010000010001100000000000",--13384
"111110001110001001110010000000000000",--13385
"111110001100001000110001100000000000",--13386
"111110001000010000110001100000000000",--13387
"010110000111000000000000000000001111",--13388
"001101001000000001000000000000000110",--13389
"011100001001000000000000000000000110",--13390
"111110000110100000000001100000000000",--13391
"111110001110010000110001100000000000",--13392
"001111001010000001000000000000000100",--13393
"111110000110001001000001100000000000",--13394
"001011000000000000110000000100101111",--13395
"000101000000000000000011010001011010",--13396
"111110000110100000000001100000000000",--13397
"111110001110000000110001100000000000",--13398
"001111001010000001000000000000000100",--13399
"111110000110001001000001100000000000",--13400
"001011000000000000110000000100101111",--13401
"101001000000000001000000000000000001",--13402
"000101000000000000000011010001011101",--13403
"101000000001111000000010000000000000",--13404
"001111000000000000110000000100101111",--13405
"010000001001000000000000000000100110",--13406
"101111001001110001001011111001001100",--13407
"101111001001100001001100110011001101",--13408
"010110001001000000110000000000100011",--13409
"101111001001110001000011110000100011",--13410
"101111001001100001001101011100001010",--13411
"111110000110000001000001100000000000",--13412
"001111000000000001000000000101100100",--13413
"111110001000001000110010000000000000",--13414
"001111000000000001010000000100101010",--13415
"111110001000000001010010000000000000",--13416
"001111000000000001010000000101100101",--13417
"111110001010001000110010100000000000",--13418
"001111000000000001100000000100101011",--13419
"111110001010000001100010100000000000",--13420
"001111000000000001100000000101100110",--13421
"111110001100001000110001100000000000",--13422
"001111000000000001100000000100101100",--13423
"111110000110000001100001100000000000",--13424
"001001111100000000101111111111111000",--13425
"101000000001111000000000100000000000",--13426
"101110001011111000001111100000000000",--13427
"101110000111111000000010100000000000",--13428
"101110001001111000000001100000000000",--13429
"101110111111111000000010000000000000",--13430
"001001111100000111111111111111110111",--13431
"101001111100010111100000000000001010",--13432
"000111000000000000000000011110001000",--13433
"101001111100000111100000000000001010",--13434
"001101111100000111111111111111110111",--13435
"011100000011000000000000000001101001",--13436
"101001000000000000010000000000000001",--13437
"001101111100000000101111111111111000",--13438
"101001111100010111100000000000001010",--13439
"000111000000000000000000100011100001",--13440
"101001111100000111100000000000001010",--13441
"001101111100000111111111111111110111",--13442
"011100000011000000000000000001100010",--13443
"000101000000000000000011010010001111",--13444
"001101000110000000110000000101101101",--13445
"001101000110000000110000000000000110",--13446
"010000000111000000000000000000000111",--13447
"101001000000000000010000000000000001",--13448
"001001111100000111111111111111111000",--13449
"101001111100010111100000000000001001",--13450
"000111000000000000000000100011100001",--13451
"101001111100000111100000000000001001",--13452
"001101111100000111111111111111111000",--13453
"011100000011000000000000000001010111",--13454
"001101111100000000011111111111111010",--13455
"001101000010000000100000000000000010",--13456
"010011000101000000000000000000001111",--13457
"001101000100000000100000000100110001",--13458
"101000000001111000000000100000000000",--13459
"001001111100000111111111111111111000",--13460
"101001111100010111100000000000001001",--13461
"000111000000000000000000100011100001",--13462
"101001111100000111100000000000001001",--13463
"001101111100000111111111111111111000",--13464
"011100000011000000000000000001001100",--13465
"101001000000000000010000000000000011",--13466
"001101111100000000101111111111111010",--13467
"101001111100010111100000000000001001",--13468
"000111000000000000000000110101111110",--13469
"101001111100000111100000000000001001",--13470
"001101111100000111111111111111111000",--13471
"011100000011000000000000000001000101",--13472
"101001000000000000010000000000000001",--13473
"001101111100000000101111111111111001",--13474
"001001111100000111111111111111111000",--13475
"101001111100010111100000000000001001",--13476
"000111000000000000000000111111111011",--13477
"101001111100000111100000000000001001",--13478
"001101111100000111111111111111111000",--13479
"011100000011000000000000000000111101",--13480
"001101111100000000011111111111111100",--13481
"001101000010000000010000000000000000",--13482
"001111000000000000110000000100100110",--13483
"001111000010000001000000000000000000",--13484
"111110000110001001000001100000000000",--13485
"001111000000000001000000000100100111",--13486
"001111000010000001010000000000000001",--13487
"111110001000001001010010000000000000",--13488
"111110000110000001000001100000000000",--13489
"001111000000000001000000000100101000",--13490
"001111000010000001010000000000000010",--13491
"111110001000001001010010000000000000",--13492
"111110000110000001000001100000000000",--13493
"001101111100000000101111111111111011",--13494
"001111000100000001000000000000000010",--13495
"001111111100000001011111111111111101",--13496
"111110001000001001010011000000000000",--13497
"111110001100001000110001100000000000",--13498
"001101111100000000101111111111111110",--13499
"001111000100000001100000000000000000",--13500
"001111000010000001110000000000000000",--13501
"111110001100001001110011000000000000",--13502
"001111000100000001110000000000000001",--13503
"001111000010000010000000000000000001",--13504
"111110001110001010000011100000000000",--13505
"111110001100000001110011000000000000",--13506
"001111000100000001110000000000000010",--13507
"001111000010000010000000000000000010",--13508
"111110001110001010000011100000000000",--13509
"111110001100000001110011000000000000",--13510
"111110001000001001100010000000000000",--13511
"010110000111000000000000000000001111",--13512
"001111000000000001100000000100011101",--13513
"001111000000000001110000000100100011",--13514
"111110000110001001110011100000000000",--13515
"111110001100000001110011000000000000",--13516
"001011000000000001100000000100011101",--13517
"001111000000000001100000000100011110",--13518
"001111000000000001110000000100100100",--13519
"111110000110001001110011100000000000",--13520
"111110001100000001110011000000000000",--13521
"001011000000000001100000000100011110",--13522
"001111000000000001100000000100011111",--13523
"001111000000000001110000000100100101",--13524
"111110000110001001110001100000000000",--13525
"111110001100000000110001100000000000",--13526
"001011000000000000110000000100011111",--13527
"010110001001000000000000000000001101",--13528
"111110001000001001000001100000000000",--13529
"111110000110001000110001100000000000",--13530
"001111111100000001001111111111111111",--13531
"111110000110001001000001100000000000",--13532
"001111000000000001100000000100011101",--13533
"111110001100000000110011000000000000",--13534
"001011000000000001100000000100011101",--13535
"001111000000000001100000000100011110",--13536
"111110001100000000110011000000000000",--13537
"001011000000000001100000000100011110",--13538
"001111000000000001100000000100011111",--13539
"111110001100000000110001100000000000",--13540
"001011000000000000110000000100011111",--13541
"001101111100000000010000000000000000",--13542
"101001000010010000010000000000000001",--13543
"010111000010000000001111100000000000",--13544
"001101000010000000100000000000000100",--13545
"001101000100000000110000000000000001",--13546
"101111000111110000110100111001101110",--13547
"101111000111100000110110101100101000",--13548
"001011000000000000110000000100101101",--13549
"001101000000000001000000000100110000",--13550
"001101001000000001010000000000000000",--13551
"001101001010000001100000000000000000",--13552
"001001111100000000011111111111111010",--13553
"001001111100000000111111111111111001",--13554
"001001111100000000101111111111111000",--13555
"010011001101000000000000000010000000",--13556
"001001111100000001001111111111110111",--13557
"011111001101011000110000000000001000",--13558
"101000001011111000000001000000000000",--13559
"101001000000000000010000000000000001",--13560
"001001111100000111111111111111110110",--13561
"101001111100010111100000000000001011",--13562
"000111000000000000000010101111001101",--13563
"101001111100000111100000000000001011",--13564
"001101111100000111111111111111110110",--13565
"000101000000000000000011010101101101",--13566
"001101001100000001110000000101101101",--13567
"001101001110000010000000000000001010",--13568
"001111010000000000110000000000000000",--13569
"001111010000000001000000000000000001",--13570
"001111010000000001010000000000000010",--13571
"001101000110000010010000000000000001",--13572
"001100010010000001100011000000000000",--13573
"001101001110000010010000000000000001",--13574
"011111010011000000010000000000111000",--13575
"001101000110000010000000000000000000",--13576
"001111001100000001100000000000000000",--13577
"111110001100010000110011000000000000",--13578
"001111001100000001110000000000000001",--13579
"111110001100001001110011000000000000",--13580
"001111010000000001110000000000000001",--13581
"111110001100001001110011100000000000",--13582
"111110001110000001000011100000000001",--13583
"001101001110000001110000000000000100",--13584
"001111001110000010000000000000000001",--13585
"010110010001000001110000000000000111",--13586
"001111010000000001110000000000000010",--13587
"111110001100001001110011100000000000",--13588
"111110001110000001010011100000000001",--13589
"001111001110000010000000000000000010",--13590
"010110010001000001110000000000000010",--13591
"001111001100000001110000000000000001",--13592
"011110001111000000000000000000100100",--13593
"001111001100000001100000000000000010",--13594
"111110001100010001000011000000000000",--13595
"001111001100000001110000000000000011",--13596
"111110001100001001110011000000000000",--13597
"001111010000000001110000000000000000",--13598
"111110001100001001110011100000000000",--13599
"111110001110000000110011100000000001",--13600
"001111001110000010000000000000000000",--13601
"010110010001000001110000000000000111",--13602
"001111010000000001110000000000000010",--13603
"111110001100001001110011100000000000",--13604
"111110001110000001010011100000000001",--13605
"001111001110000010000000000000000010",--13606
"010110010001000001110000000000000010",--13607
"001111001100000001110000000000000011",--13608
"011110001111000000000000000000010010",--13609
"001111001100000001100000000000000100",--13610
"111110001100010001010010100000000000",--13611
"001111001100000001100000000000000101",--13612
"111110001010001001100010100000000000",--13613
"001111010000000001100000000000000000",--13614
"111110001010001001100011000000000000",--13615
"111110001100000000110001100000000001",--13616
"001111001110000001100000000000000000",--13617
"010110001101000000110000000000111010",--13618
"001111010000000000110000000000000001",--13619
"111110001010001000110001100000000000",--13620
"111110000110000001000001100000000001",--13621
"001111001110000001000000000000000001",--13622
"010110001001000000110000000000110101",--13623
"001111001100000000110000000000000101",--13624
"010010000111000000000000000000110011",--13625
"001011000000000001010000000100101111",--13626
"000101000000000000000011010101100011",--13627
"001011000000000001100000000100101111",--13628
"000101000000000000000011010101100011",--13629
"001011000000000001100000000100101111",--13630
"000101000000000000000011010101100011",--13631
"011111010011000000100000000000000110",--13632
"001111001100000000110000000000000000",--13633
"011010000111000000000000000000101010",--13634
"001111010000000001000000000000000011",--13635
"111110000110001001000001100000000000",--13636
"001011000000000000110000000100101111",--13637
"000101000000000000000011010101100011",--13638
"001111001100000001100000000000000000",--13639
"010010001101000000000000000000100100",--13640
"001111001100000001110000000000000001",--13641
"111110001110001000110001100000000000",--13642
"001111001100000001110000000000000010",--13643
"111110001110001001000010000000000000",--13644
"111110000110000001000001100000000000",--13645
"001111001100000001000000000000000011",--13646
"111110001000001001010010000000000000",--13647
"111110000110000001000001100000000000",--13648
"001111010000000001000000000000000011",--13649
"111110000110001000110010100000000000",--13650
"111110001100001001000010000000000000",--13651
"111110001010010001000010000000000000",--13652
"010110001001000000000000000000010111",--13653
"001101001110000001110000000000000110",--13654
"011100001111000000000000000000000110",--13655
"111110001000100000000010000000000000",--13656
"111110000110010001000001100000000000",--13657
"001111001100000001000000000000000100",--13658
"111110000110001001000001100000000000",--13659
"001011000000000000110000000100101111",--13660
"000101000000000000000011010101100011",--13661
"111110001000100000000010000000000000",--13662
"111110000110000001000001100000000000",--13663
"001111001100000001000000000000000100",--13664
"111110000110001001000001100000000000",--13665
"001011000000000000110000000100101111",--13666
"001111000000000000110000000100101111",--13667
"001111000000000001000000000100101101",--13668
"010110001001000000110000000000000111",--13669
"101000001011111000000001000000000000",--13670
"101001000000000000010000000000000001",--13671
"001001111100000111111111111111110110",--13672
"101001111100010111100000000000001011",--13673
"000111000000000000000010101111001101",--13674
"101001111100000111100000000000001011",--13675
"001101111100000111111111111111110110",--13676
"101001000000000000010000000000000001",--13677
"001101111100000000101111111111110111",--13678
"001101111100000000111111111111111001",--13679
"001001111100000111111111111111110110",--13680
"101001111100010111100000000000001011",--13681
"000111000000000000000010110111111111",--13682
"101001111100000111100000000000001011",--13683
"001101111100000111111111111111110110",--13684
"001111000000000000110000000100101101",--13685
"101111001001110001001011110111001100",--13686
"101111001001100001001100110011001101",--13687
"010110000111000001000000000001001111",--13688
"101111001001110001000100110010111110",--13689
"101111001001100001001011110000100000",--13690
"010110001001000000110000000001001100",--13691
"001101000000000000010000000100101001",--13692
"101000000011000000010000100010000010",--13693
"001101000000000000100000000100101110",--13694
"101000000010000000100000100000000000",--13695
"001101111100000000101111111111111000",--13696
"001101000100000000110000000000000000",--13697
"011100000011000000110000000001000101",--13698
"101000000001111000000000100000000000",--13699
"001101000000000000100000000100110000",--13700
"001001111100000111111111111111110111",--13701
"101001111100010111100000000000001010",--13702
"000111000000000000000000111111111011",--13703
"101001111100000111100000000000001010",--13704
"001101111100000111111111111111110111",--13705
"011100000011000000000000000000111101",--13706
"001101111100000000011111111111111001",--13707
"001101000010000000010000000000000000",--13708
"001111000000000000110000000100100110",--13709
"001111000010000001000000000000000000",--13710
"111110000110001001000001100000000000",--13711
"001111000000000001000000000100100111",--13712
"001111000010000001010000000000000001",--13713
"111110001000001001010010000000000000",--13714
"111110000110000001000001100000000000",--13715
"001111000000000001000000000100101000",--13716
"001111000010000001010000000000000010",--13717
"111110001000001001010010000000000000",--13718
"111110000110000001000001100000000000",--13719
"001101111100000000101111111111111000",--13720
"001111000100000001000000000000000010",--13721
"001111111100000001011111111111111101",--13722
"111110001000001001010011000000000000",--13723
"111110001100001000110001100000000000",--13724
"001101111100000000101111111111111110",--13725
"001111000100000001100000000000000000",--13726
"001111000010000001110000000000000000",--13727
"111110001100001001110011000000000000",--13728
"001111000100000001110000000000000001",--13729
"001111000010000010000000000000000001",--13730
"111110001110001010000011100000000000",--13731
"111110001100000001110011000000000000",--13732
"001111000100000001110000000000000010",--13733
"001111000010000010000000000000000010",--13734
"111110001110001010000011100000000000",--13735
"111110001100000001110011000000000000",--13736
"111110001000001001100010000000000000",--13737
"010110000111000000000000000000001111",--13738
"001111000000000001100000000100011101",--13739
"001111000000000001110000000100100011",--13740
"111110000110001001110011100000000000",--13741
"111110001100000001110011000000000000",--13742
"001011000000000001100000000100011101",--13743
"001111000000000001100000000100011110",--13744
"001111000000000001110000000100100100",--13745
"111110000110001001110011100000000000",--13746
"111110001100000001110011000000000000",--13747
"001011000000000001100000000100011110",--13748
"001111000000000001100000000100011111",--13749
"001111000000000001110000000100100101",--13750
"111110000110001001110001100000000000",--13751
"111110001100000000110001100000000000",--13752
"001011000000000000110000000100011111",--13753
"010110001001000000000000000000001101",--13754
"111110001000001001000001100000000000",--13755
"111110000110001000110001100000000000",--13756
"001111111100000001001111111111111111",--13757
"111110000110001001000001100000000000",--13758
"001111000000000001100000000100011101",--13759
"111110001100000000110011000000000000",--13760
"001011000000000001100000000100011101",--13761
"001111000000000001100000000100011110",--13762
"111110001100000000110011000000000000",--13763
"001011000000000001100000000100011110",--13764
"001111000000000001100000000100011111",--13765
"111110001100000000110001100000000000",--13766
"001011000000000000110000000100011111",--13767
"001101111100000000011111111111111010",--13768
"101001000010010000010000000000000001",--13769
"001111111100000000111111111111111101",--13770
"001111111100000001001111111111111111",--13771
"001101111100000000101111111111111110",--13772
"010111000010000000001111100000000000",--13773
"000101000000000000000011001000010101",--13774
"011011000010000001011111100000000000",--13775
"001101000110000001000000000000000010",--13776
"101111001011110001010100111001101110",--13777
"101111001011100001010110101100101000",--13778
"001011000000000001010000000100101101",--13779
"001101000000000001100000000100110000",--13780
"001011111100000001000000000000000000",--13781
"001001111100000000111111111111111111",--13782
"001011111100000000111111111111111110",--13783
"001001111100000000101111111111111101",--13784
"001001111100000001001111111111111100",--13785
"001001111100000000011111111111111011",--13786
"101000000101111000000001100000000000",--13787
"101000000001111000000000100000000000",--13788
"101000001101111000000001000000000000",--13789
"001001111100000111111111111111111010",--13790
"101001111100010111100000000000000111",--13791
"000111000000000000000010000001010110",--13792
"101001111100000111100000000000000111",--13793
"001101111100000111111111111111111010",--13794
"001111000000000000110000000100101101",--13795
"101111001001110001001011110111001100",--13796
"101111001001100001001100110011001101",--13797
"010110000111000001000000000000010110",--13798
"101111001001110001000100110010111110",--13799
"101111001001100001001011110000100000",--13800
"010110001001000000110000000000010011",--13801
"001101000000000000010000000100101001",--13802
"001101000010000000100000000101101101",--13803
"001101000100000000110000000000000111",--13804
"001111000110000000110000000000000000",--13805
"001111111100000001001111111111111110",--13806
"111110000110001001000001100000000000",--13807
"001101000100000001000000000000000001",--13808
"011111001001000000010000000000110100",--13809
"001101000000000001000000000100101110",--13810
"001011000000000000000000000100100110",--13811
"001011000000000000000000000100100111",--13812
"001011000000000000000000000100101000",--13813
"101001001000010001010000000000000001",--13814
"101001001000010001000000000000000001",--13815
"001101111100000001101111111111111101",--13816
"001110001100000001000010100000000000",--13817
"011110001011000000000000000000100100",--13818
"101110000001111000000010100000000000",--13819
"000101000000000000000011011000100011",--13820
"101001000000000000011111111111111111",--13821
"001101111100000000101111111111111011",--13822
"001101111100000001001111111111111100",--13823
"001000001000000000100000100000000000",--13824
"010000000100000000001111100000000000",--13825
"001101111100000000011111111111111101",--13826
"001111000010000000110000000000000000",--13827
"001111000000000001000000000101100100",--13828
"111110000110001001000001100000000000",--13829
"001111000010000001000000000000000001",--13830
"001111000000000001010000000101100101",--13831
"111110001000001001010010000000000000",--13832
"111110000110000001000001100000000000",--13833
"001111000010000001000000000000000010",--13834
"001111000000000001010000000101100110",--13835
"111110001000001001010010000000000000",--13836
"111110000110000001000001100000000010",--13837
"010110000110000000001111100000000000",--13838
"111110000110001000110010000000000000",--13839
"111110001000001000110001100000000000",--13840
"001111111100000001001111111111111110",--13841
"111110000110001001000001100000000000",--13842
"001111000000000001000000000101100011",--13843
"111110000110001001000001100000000000",--13844
"001111000000000001000000000100011101",--13845
"111110001000000000110010000000000000",--13846
"001011000000000001000000000100011101",--13847
"001111000000000001000000000100011110",--13848
"111110001000000000110010000000000000",--13849
"001011000000000001000000000100011110",--13850
"001111000000000001000000000100011111",--13851
"111110001000000000110001100000000000",--13852
"001011000000000000110000000100011111",--13853
"000100000000000000001111100000000000",--13854
"010110001011000000000000000000000010",--13855
"101110000011111000000010100000000000",--13856
"000101000000000000000011011000100011",--13857
"101110000101111000000010100000000000",--13858
"101110001011111000000010100000000010",--13859
"001011001010000001010000000100100110",--13860
"000101000000000000000011011001111100",--13861
"011111001001000000100000000000001000",--13862
"001101000100000001000000000000000100",--13863
"001111001000010001010000000000000000",--13864
"001011000000000001010000000100100110",--13865
"001111001000010001010000000000000001",--13866
"001011000000000001010000000100100111",--13867
"001111001000010001010000000000000010",--13868
"001011000000000001010000000100101000",--13869
"000101000000000000000011011001111100",--13870
"001111000000000001010000000100101010",--13871
"001101000100000001000000000000000101",--13872
"001111001000000001100000000000000000",--13873
"111110001010010001100010100000000000",--13874
"001111000000000001100000000100101011",--13875
"001111001000000001110000000000000001",--13876
"111110001100010001110011000000000000",--13877
"001111000000000001110000000100101100",--13878
"001111001000000010000000000000000010",--13879
"111110001110010010000011100000000000",--13880
"001101000100000001000000000000000100",--13881
"001111001000000010000000000000000000",--13882
"111110001010001010000100000000000000",--13883
"001111001000000010010000000000000001",--13884
"111110001100001010010100100000000000",--13885
"001111001000000010100000000000000010",--13886
"111110001110001010100101000000000000",--13887
"001101000100000001000000000000000011",--13888
"011100001001000000000000000000000100",--13889
"001011000000000010000000000100100110",--13890
"001011000000000010010000000100100111",--13891
"001011000000000010100000000100101000",--13892
"000101000000000000000011011001100010",--13893
"001101000100000001000000000000001001",--13894
"001111001000000010110000000000000010",--13895
"111110001100001010110101100000000000",--13896
"001111001000000011000000000000000001",--13897
"111110001110001011000110000000000000",--13898
"111110010110000011000101100000000000",--13899
"101111000001110011000011111100000000",--13900
"111110010110001011000101100000000000",--13901
"111110010000000010110100000000000000",--13902
"001011000000000010000000000100100110",--13903
"001111001000000010000000000000000010",--13904
"111110001010001010000100000000000000",--13905
"001111001000000010110000000000000000",--13906
"111110001110001010110011100000000000",--13907
"111110010000000001110011100000000000",--13908
"101111000001110010000011111100000000",--13909
"111110001110001010000011100000000000",--13910
"111110010010000001110011100000000000",--13911
"001011000000000001110000000100100111",--13912
"001111001000000001110000000000000001",--13913
"111110001010001001110010100000000000",--13914
"001111001000000001110000000000000000",--13915
"111110001100001001110011000000000000",--13916
"111110001010000001100010100000000000",--13917
"101111000001110001100011111100000000",--13918
"111110001010001001100010100000000000",--13919
"111110010100000001010010100000000000",--13920
"001011000000000001010000000100101000",--13921
"001111000000000001010000000100100110",--13922
"111110001010001001010010100000000000",--13923
"001111000000000001100000000100100111",--13924
"111110001100001001100011000000000000",--13925
"111110001010000001100010100000000000",--13926
"001111000000000001100000000100101000",--13927
"111110001100001001100011000000000000",--13928
"111110001010000001100010100000000000",--13929
"111110001010100000000010100000000000",--13930
"011110001011000000000000000000000010",--13931
"101110000011111000000010100000000000",--13932
"000101000000000000000011011001110011",--13933
"001101000100000001000000000000000110",--13934
"011100001001000000000000000000000010",--13935
"111110001010011000000010100000000000",--13936
"000101000000000000000011011001110011",--13937
"111110001010011000000010100000000010",--13938
"001111000000000001100000000100100110",--13939
"111110001100001001010011000000000000",--13940
"001011000000000001100000000100100110",--13941
"001111000000000001100000000100100111",--13942
"111110001100001001010011000000000000",--13943
"001011000000000001100000000100100111",--13944
"001111000000000001100000000100101000",--13945
"111110001100001001010010100000000000",--13946
"001011000000000001010000000100101000",--13947
"001111000000000001010000000100101010",--13948
"001011000000000001010000000100010101",--13949
"001111000000000001010000000100101011",--13950
"001011000000000001010000000100010110",--13951
"001111000000000001010000000100101100",--13952
"001011000000000001010000000100010111",--13953
"001101000100000001000000000000000000",--13954
"001101000100000001010000000000001000",--13955
"001111001010000001010000000000000000",--13956
"001011000000000001010000000100100011",--13957
"001111001010000001010000000000000001",--13958
"001011000000000001010000000100100100",--13959
"001111001010000001010000000000000010",--13960
"001011000000000001010000000100100101",--13961
"001001111100000000101111111111111010",--13962
"001011111100000000111111111111111001",--13963
"001001111100000000111111111111111000",--13964
"001001111100000000011111111111110111",--13965
"011111001001000000010000000000100011",--13966
"001111000000000001010000000100101010",--13967
"001101000100000001000000000000000101",--13968
"001111001000000001100000000000000000",--13969
"111110001010010001100010100000000000",--13970
"101111001101110001100011110101001100",--13971
"101111001101100001101100110011001101",--13972
"111110001010001001100011000000000000",--13973
"101110001100110000000011000000000000",--13974
"101111000001110001110100000110100000",--13975
"111110001100001001110011000000000000",--13976
"111110001010010001100010100000000000",--13977
"101111000001110001100100000100100000",--13978
"001111000000000001110000000100101100",--13979
"001111001000000010000000000000000010",--13980
"111110001110010010000011100000000000",--13981
"101111010001110010000011110101001100",--13982
"101111010001100010001100110011001101",--13983
"111110001110001010000100000000000000",--13984
"101110010000110000000100000000000000",--13985
"101111000001110010010100000110100000",--13986
"111110010000001010010100000000000000",--13987
"111110001110010010000011100000000000",--13988
"101111000001110010000100000100100000",--13989
"010110001101000001010000000000000101",--13990
"010110010001000001110000000000000010",--13991
"101111000001110001010100001101111111",--13992
"000101000000000000000011011010110000",--13993
"101110000001111000000010100000000000",--13994
"000101000000000000000011011010110000",--13995
"010110010001000001110000000000000010",--13996
"101110000001111000000010100000000000",--13997
"000101000000000000000011011010110000",--13998
"101111000001110001010100001101111111",--13999
"001011000000000001010000000100100100",--14000
"000101000000000000000011011111010110",--14001
"011111001001000000100000000000010000",--14002
"001111000000000001010000000100101011",--14003
"101111000001110001100011111010000000",--14004
"111110001010001001100010100000000000",--14005
"101110001011111000000001100000000000",--14006
"001001111100000111111111111111110110",--14007
"000111000000000000000111011000000010",--14008
"001101111100000111111111111111110110",--14009
"111110000110001000110001100000000000",--14010
"101111000001110001000100001101111111",--14011
"111110001000001000110010000000000000",--14012
"001011000000000001000000000100100011",--14013
"101111000001110001000100001101111111",--14014
"111110000110010000010001100000000010",--14015
"111110001000001000110001100000000000",--14016
"001011000000000000110000000100100100",--14017
"000101000000000000000011011111010110",--14018
"011111001001000000110000000000100000",--14019
"001111000000000001010000000100101010",--14020
"001101000100000001000000000000000101",--14021
"001111001000000001100000000000000000",--14022
"111110001010010001100010100000000000",--14023
"001111000000000001100000000100101100",--14024
"001111001000000001110000000000000010",--14025
"111110001100010001110011000000000000",--14026
"111110001010001001010010100000000000",--14027
"111110001100001001100011000000000000",--14028
"111110001010000001100010100000000000",--14029
"111110001010100000000010100000000000",--14030
"101111001101110001100011110111001100",--14031
"101111001101100001101100110011001100",--14032
"111110001010001001100010100000000000",--14033
"101110001010110000000011000000000000",--14034
"111110001010010001100010100000000000",--14035
"101111001101110001100100000001001001",--14036
"101111001101100001100000111111011011",--14037
"111110001010001001100010100000000000",--14038
"101110001011111000000001100000000000",--14039
"001001111100000111111111111111110110",--14040
"000111000000000000000111010110111000",--14041
"001101111100000111111111111111110110",--14042
"111110000110001000110001100000000000",--14043
"101111000001110001000100001101111111",--14044
"111110000110001001000010000000000000",--14045
"001011000000000001000000000100100100",--14046
"111110000110010000010001100000000010",--14047
"101111000001110001000100001101111111",--14048
"111110000110001001000001100000000000",--14049
"001011000000000000110000000100100101",--14050
"000101000000000000000011011111010110",--14051
"011111001001000001000000000011110001",--14052
"001111000000000001010000000100101010",--14053
"001101000100000001000000000000000101",--14054
"001111001000000001100000000000000000",--14055
"111110001010010001100010100000000000",--14056
"001101000100000001010000000000000100",--14057
"001111001010000001100000000000000000",--14058
"111110001100100000000011000000000000",--14059
"111110001010001001100010100000000000",--14060
"001111000000000001100000000100101100",--14061
"001111001000000001110000000000000010",--14062
"111110001100010001110011000000000000",--14063
"001111001010000001110000000000000010",--14064
"111110001110100000000011100000000000",--14065
"111110001100001001110011000000000000",--14066
"111110001010001001010011100000000000",--14067
"111110001100001001100100000000000000",--14068
"111110001110000010000011100000000000",--14069
"101110001011111000000100000000000001",--14070
"101111010011110010010011100011010001",--14071
"101111010011100010011011011100010111",--14072
"010110010011000010000000000000000010",--14073
"101111000001110001010100000101110000",--14074
"000101000000000000000011011101011000",--14075
"111110001010011000000010100000000000",--14076
"111110001100001001010010100000000001",--14077
"010110001011000000010000000000000010",--14078
"101001000000000001100000000000000001",--14079
"000101000000000000000011011100000110",--14080
"011010001011000000100000000000000010",--14081
"101001000000000001101111111111111111",--14082
"000101000000000000000011011100000110",--14083
"101000000001111000000011000000000000",--14084
"000101000000000000000011011100000111",--14085
"111110001010011000000010100000000000",--14086
"111110001010001001010011000000000000",--14087
"101111000001110010000100001011110010",--14088
"111110010000001001100100000000000000",--14089
"101111010011110010010011110100110010",--14090
"101111010011100010010001011001000011",--14091
"111110010000001010010100000000000000",--14092
"101111000001110010010100001011001000",--14093
"111110010010001001100100100000000000",--14094
"101111000001110010100100000110101000",--14095
"111110010100000010000100000000000000",--14096
"111110010000011000000100000000000000",--14097
"111110010010001010000100000000000000",--14098
"101111000001110010010100001010100010",--14099
"111110010010001001100100100000000000",--14100
"101111000001110010100100000110011000",--14101
"111110010100000010000100000000000000",--14102
"111110010000011000000100000000000000",--14103
"111110010010001010000100000000000000",--14104
"101111000001110010010100001010000000",--14105
"111110010010001001100100100000000000",--14106
"101111000001110010100100000110001000",--14107
"111110010100000010000100000000000000",--14108
"111110010000011000000100000000000000",--14109
"111110010010001010000100000000000000",--14110
"101111000001110010010100001001000100",--14111
"111110010010001001100100100000000000",--14112
"101111000001110010100100000101110000",--14113
"111110010100000010000100000000000000",--14114
"111110010000011000000100000000000000",--14115
"111110010010001010000100000000000000",--14116
"101111000001110010010100001000010000",--14117
"111110010010001001100100100000000000",--14118
"101111000001110010100100000101010000",--14119
"111110010100000010000100000000000000",--14120
"111110010000011000000100000000000000",--14121
"111110010010001010000100000000000000",--14122
"101111000001110010010100000111001000",--14123
"111110010010001001100100100000000000",--14124
"101111000001110010100100000100110000",--14125
"111110010100000010000100000000000000",--14126
"111110010000011000000100000000000000",--14127
"111110010010001010000100000000000000",--14128
"101111000001110010010100000110000000",--14129
"111110010010001001100100100000000000",--14130
"101111000001110010100100000100010000",--14131
"111110010100000010000100000000000000",--14132
"111110010000011000000100000000000000",--14133
"111110010010001010000100000000000000",--14134
"101111000001110010010100000100010000",--14135
"111110010010001001100100100000000000",--14136
"101111000001110010100100000011100000",--14137
"111110010100000010000100000000000000",--14138
"111110010000011000000100000000000000",--14139
"111110010010001010000100000000000000",--14140
"101111000001110010010100000010000000",--14141
"111110010010001001100100100000000000",--14142
"101111000001110010100100000010100000",--14143
"111110010100000010000100000000000000",--14144
"111110010000011000000100000000000000",--14145
"111110010010001010000100000000000000",--14146
"101111000001110010010100000001000000",--14147
"111110010010000010000100000000000000",--14148
"111110010000011000000100000000000000",--14149
"111110001100001010000011000000000000",--14150
"111110001100000000010011000000000000",--14151
"111110001100011000000011000000000000",--14152
"111110001010001001100010100000000000",--14153
"010100001101000000000000000000000100",--14154
"101111001101110001100011111111001001",--14155
"101111001101100001100000111111011010",--14156
"111110001100010001010010100000000000",--14157
"000101000000000000000011011101010011",--14158
"011000001101000000000000000000000011",--14159
"101111001101110001101011111111001001",--14160
"101111001101100001100000111111011010",--14161
"111110001100010001010010100000000000",--14162
"101111000001110001100100000111110000",--14163
"111110001010001001100010100000000000",--14164
"101111001101110001100011111010100010",--14165
"101111001101100001101111100110000010",--14166
"111110001010001001100010100000000000",--14167
"101110001010110000000011000000000000",--14168
"111110001010010001100010100000000000",--14169
"101110001111111000000011000000000001",--14170
"101111010001110010000011100011010001",--14171
"101111010001100010001011011100010111",--14172
"010110010001000001100000000000000010",--14173
"101111000001110001100100000101110000",--14174
"000101000000000000000011011111000010",--14175
"001111000000000001100000000100101011",--14176
"001111001000000010000000000000000001",--14177
"111110001100010010000011000000000000",--14178
"001111001010000010000000000000000001",--14179
"111110010000100000000100000000000000",--14180
"111110001100001010000011000000000000",--14181
"111110001110011000000011100000000000",--14182
"111110001100001001110011000000000001",--14183
"010110001101000000010000000000000010",--14184
"101001000000000001000000000000000001",--14185
"000101000000000000000011011101110000",--14186
"011010001101000000100000000000000010",--14187
"101001000000000001001111111111111111",--14188
"000101000000000000000011011101110000",--14189
"101000000001111000000010000000000000",--14190
"000101000000000000000011011101110001",--14191
"111110001100011000000011000000000000",--14192
"111110001100001001100011100000000000",--14193
"101111000001110010000100001011110010",--14194
"111110010000001001110100000000000000",--14195
"101111010011110010010011110100110010",--14196
"101111010011100010010001011001000011",--14197
"111110010000001010010100000000000000",--14198
"101111000001110010010100001011001000",--14199
"111110010010001001110100100000000000",--14200
"101111000001110010100100000110101000",--14201
"111110010100000010000100000000000000",--14202
"111110010000011000000100000000000000",--14203
"111110010010001010000100000000000000",--14204
"101111000001110010010100001010100010",--14205
"111110010010001001110100100000000000",--14206
"101111000001110010100100000110011000",--14207
"111110010100000010000100000000000000",--14208
"111110010000011000000100000000000000",--14209
"111110010010001010000100000000000000",--14210
"101111000001110010010100001010000000",--14211
"111110010010001001110100100000000000",--14212
"101111000001110010100100000110001000",--14213
"111110010100000010000100000000000000",--14214
"111110010000011000000100000000000000",--14215
"111110010010001010000100000000000000",--14216
"101111000001110010010100001001000100",--14217
"111110010010001001110100100000000000",--14218
"101111000001110010100100000101110000",--14219
"111110010100000010000100000000000000",--14220
"111110010000011000000100000000000000",--14221
"111110010010001010000100000000000000",--14222
"101111000001110010010100001000010000",--14223
"111110010010001001110100100000000000",--14224
"101111000001110010100100000101010000",--14225
"111110010100000010000100000000000000",--14226
"111110010000011000000100000000000000",--14227
"111110010010001010000100000000000000",--14228
"101111000001110010010100000111001000",--14229
"111110010010001001110100100000000000",--14230
"101111000001110010100100000100110000",--14231
"111110010100000010000100000000000000",--14232
"111110010000011000000100000000000000",--14233
"111110010010001010000100000000000000",--14234
"101111000001110010010100000110000000",--14235
"111110010010001001110100100000000000",--14236
"101111000001110010100100000100010000",--14237
"111110010100000010000100000000000000",--14238
"111110010000011000000100000000000000",--14239
"111110010010001010000100000000000000",--14240
"101111000001110010010100000100010000",--14241
"111110010010001001110100100000000000",--14242
"101111000001110010100100000011100000",--14243
"111110010100000010000100000000000000",--14244
"111110010000011000000100000000000000",--14245
"111110010010001010000100000000000000",--14246
"101111000001110010010100000010000000",--14247
"111110010010001001110100100000000000",--14248
"101111000001110010100100000010100000",--14249
"111110010100000010000100000000000000",--14250
"111110010000011000000100000000000000",--14251
"111110010010001010000100000000000000",--14252
"101111000001110010010100000001000000",--14253
"111110010010000010000100000000000000",--14254
"111110010000011000000100000000000000",--14255
"111110001110001010000011100000000000",--14256
"111110001110000000010011100000000000",--14257
"111110001110011000000011100000000000",--14258
"111110001100001001110011000000000000",--14259
"010100001001000000000000000000000100",--14260
"101111001111110001110011111111001001",--14261
"101111001111100001110000111111011010",--14262
"111110001110010001100011000000000000",--14263
"000101000000000000000011011110111101",--14264
"011000001001000000000000000000000011",--14265
"101111001111110001111011111111001001",--14266
"101111001111100001110000111111011010",--14267
"111110001110010001100011000000000000",--14268
"101111000001110001110100000111110000",--14269
"111110001100001001110011000000000000",--14270
"101111001111110001110011111010100010",--14271
"101111001111100001111111100110000010",--14272
"111110001100001001110011000000000000",--14273
"101110001100110000000011100000000000",--14274
"111110001100010001110011000000000000",--14275
"101111001111110001110011111000011001",--14276
"101111001111100001111001100110011010",--14277
"101111000001110010000011111100000000",--14278
"111110010000010001010010100000000000",--14279
"111110001010001001010010100000000000",--14280
"111110001110010001010010100000000000",--14281
"101111000001110001110011111100000000",--14282
"111110001110010001100011000000000000",--14283
"111110001100001001100011000000000000",--14284
"111110001010010001100010100000000000",--14285
"011010001011000000000000000000000001",--14286
"101110000001111000000010100000000000",--14287
"101111000001110001100100001101111111",--14288
"111110001100001001010010100000000000",--14289
"101111001101110001100100000001010101",--14290
"101111001101100001100101010101010101",--14291
"111110001010001001100010100000000000",--14292
"001011000000000001010000000100100101",--14293
"001101111100000000011111111111110111",--14294
"101000000011000000010000100010000010",--14295
"001101000000000000100000000100101110",--14296
"101000000010000000100000100000000000",--14297
"001101111100000000101111111111111011",--14298
"001101111100000001001111111111111100",--14299
"001000001000000000100000100000000000",--14300
"001101111100000000111111111111111111",--14301
"001101000110000000010000000000000001",--14302
"001100000010000000100000100000000000",--14303
"001111000000000000110000000100101010",--14304
"001011000010000000110000000000000000",--14305
"001111000000000000110000000100101011",--14306
"001011000010000000110000000000000001",--14307
"001111000000000000110000000100101100",--14308
"001011000010000000110000000000000010",--14309
"001101000110000000010000000000000011",--14310
"001101111100000001011111111111111000",--14311
"001111001010000000110000000000000000",--14312
"101111000001110001000011111100000000",--14313
"010110001001000000110000000000000010",--14314
"001000000010000000100000000000000000",--14315
"000101000000000000000011100000001101",--14316
"101001000000000001100000000000000001",--14317
"001000000010000000100011000000000000",--14318
"001101000110000000010000000000000100",--14319
"001100000010000000100011000000000000",--14320
"001111000000000000110000000100100011",--14321
"001011001100000000110000000000000000",--14322
"001111000000000000110000000100100100",--14323
"001011001100000000110000000000000001",--14324
"001111000000000000110000000100100101",--14325
"001011001100000000110000000000000010",--14326
"001100000010000000100000100000000000",--14327
"101111000111110000110011101101111111",--14328
"101111000111100000111111111111111111",--14329
"001111111100000001001111111111111001",--14330
"111110000110001001000001100000000000",--14331
"001111000010000001010000000000000000",--14332
"111110001010001000110010100000000000",--14333
"001011000010000001010000000000000000",--14334
"001111000010000001010000000000000001",--14335
"111110001010001000110010100000000000",--14336
"001011000010000001010000000000000001",--14337
"001111000010000001010000000000000010",--14338
"111110001010001000110001100000000000",--14339
"001011000010000000110000000000000010",--14340
"001101000110000000010000000000000111",--14341
"001100000010000000100000100000000000",--14342
"001111000000000000110000000100100110",--14343
"001011000010000000110000000000000000",--14344
"001111000000000000110000000100100111",--14345
"001011000010000000110000000000000001",--14346
"001111000000000000110000000100101000",--14347
"001011000010000000110000000000000010",--14348
"101111000001110000111100000000000000",--14349
"001101111100000000011111111111111101",--14350
"001111000010000001000000000000000000",--14351
"001111000000000001010000000100100110",--14352
"111110001000001001010010000000000000",--14353
"001111000010000001010000000000000001",--14354
"001111000000000001100000000100100111",--14355
"111110001010001001100010100000000000",--14356
"111110001000000001010010000000000000",--14357
"001111000010000001010000000000000010",--14358
"001111000000000001100000000100101000",--14359
"111110001010001001100010100000000000",--14360
"111110001000000001010010000000000000",--14361
"111110000110001001000001100000000000",--14362
"001111000010000001000000000000000000",--14363
"001111000000000001010000000100100110",--14364
"111110000110001001010010100000000000",--14365
"111110001000000001010010000000000000",--14366
"001011000010000001000000000000000000",--14367
"001111000010000001000000000000000001",--14368
"001111000000000001010000000100100111",--14369
"111110000110001001010010100000000000",--14370
"111110001000000001010010000000000000",--14371
"001011000010000001000000000000000001",--14372
"001111000010000001000000000000000010",--14373
"001111000000000001010000000100101000",--14374
"111110000110001001010001100000000000",--14375
"111110001000000000110001100000000000",--14376
"001011000010000000110000000000000010",--14377
"001111001010000000110000000000000001",--14378
"001111111100000001001111111111111110",--14379
"111110001000001000110001100000000000",--14380
"001101000000000001100000000100110000",--14381
"001101001100000001110000000000000000",--14382
"001101001110000010000000000000000000",--14383
"001011111100000000111111111111110110",--14384
"010011010001000000000000001001101100",--14385
"001001111100000001111111111111110101",--14386
"001001111100000001101111111111110100",--14387
"010011010001011000110000000101111101",--14388
"001101010000000010010000000101101101",--14389
"001111000000000001010000000100101010",--14390
"001101010010000010100000000000000101",--14391
"001111010100000001100000000000000000",--14392
"111110001010010001100010100000000000",--14393
"001111000000000001100000000100101011",--14394
"001111010100000001110000000000000001",--14395
"111110001100010001110011000000000000",--14396
"001111000000000001110000000100101100",--14397
"001111010100000010000000000000000010",--14398
"111110001110010010000011100000000000",--14399
"001101010000000010000000000010111110",--14400
"001101010010000010100000000000000001",--14401
"011111010101000000010000000000110111",--14402
"001111010000000010000000000000000000",--14403
"111110010000010001010100000000000000",--14404
"001111010000000010010000000000000001",--14405
"111110010000001010010100000000000000",--14406
"001111000000000010010000000011111011",--14407
"111110010000001010010100100000000000",--14408
"111110010010000001100100100000000001",--14409
"001101010010000010010000000000000100",--14410
"001111010010000010100000000000000001",--14411
"010110010101000010010000000000000111",--14412
"001111000000000010010000000011111100",--14413
"111110010000001010010100100000000000",--14414
"111110010010000001110100100000000001",--14415
"001111010010000010100000000000000010",--14416
"010110010101000010010000000000000010",--14417
"001111010000000010010000000000000001",--14418
"011110010011000000000000000000100100",--14419
"001111010000000010000000000000000010",--14420
"111110010000010001100100000000000000",--14421
"001111010000000010010000000000000011",--14422
"111110010000001010010100000000000000",--14423
"001111000000000010010000000011111010",--14424
"111110010000001010010100100000000000",--14425
"111110010010000001010100100000000001",--14426
"001111010010000010100000000000000000",--14427
"010110010101000010010000000000000111",--14428
"001111000000000010010000000011111100",--14429
"111110010000001010010100100000000000",--14430
"111110010010000001110100100000000001",--14431
"001111010010000010100000000000000010",--14432
"010110010101000010010000000000000010",--14433
"001111010000000010010000000000000011",--14434
"011110010011000000000000000000010010",--14435
"001111010000000010000000000000000100",--14436
"111110010000010001110011100000000000",--14437
"001111010000000010000000000000000101",--14438
"111110001110001010000011100000000000",--14439
"001111000000000010000000000011111010",--14440
"111110001110001010000100000000000000",--14441
"111110010000000001010010100000000001",--14442
"001111010010000010000000000000000000",--14443
"010110010001000001010000000100111100",--14444
"001111000000000001010000000011111011",--14445
"111110001110001001010010100000000000",--14446
"111110001010000001100010100000000001",--14447
"001111010010000001100000000000000001",--14448
"010110001101000001010000000100110111",--14449
"001111010000000001010000000000000101",--14450
"010010001011000000000000000100110101",--14451
"001011000000000001110000000100101111",--14452
"000101000000000000000011100011000010",--14453
"001011000000000010000000000100101111",--14454
"000101000000000000000011100011000010",--14455
"001011000000000010000000000100101111",--14456
"000101000000000000000011100011000010",--14457
"011111010101000000100000000000001100",--14458
"001111010000000010000000000000000000",--14459
"011010010001000000000000000100101100",--14460
"001111010000000010000000000000000001",--14461
"111110010000001001010010100000000000",--14462
"001111010000000010000000000000000010",--14463
"111110010000001001100011000000000000",--14464
"111110001010000001100010100000000000",--14465
"001111010000000001100000000000000011",--14466
"111110001100001001110011000000000000",--14467
"111110001010000001100010100000000000",--14468
"001011000000000001010000000100101111",--14469
"000101000000000000000011100011000010",--14470
"001111010000000010000000000000000000",--14471
"010010010001000000000000000100100000",--14472
"001111010000000010010000000000000001",--14473
"111110010010001001010100100000000000",--14474
"001111010000000010100000000000000010",--14475
"111110010100001001100101000000000000",--14476
"111110010010000010100100100000000000",--14477
"001111010000000010100000000000000011",--14478
"111110010100001001110101000000000000",--14479
"111110010010000010100100100000000000",--14480
"111110001010001001010101000000000000",--14481
"001101010010000010110000000000000100",--14482
"001111010110000010110000000000000000",--14483
"111110010100001010110101000000000000",--14484
"111110001100001001100101100000000000",--14485
"001111010110000011000000000000000001",--14486
"111110010110001011000101100000000000",--14487
"111110010100000010110101000000000000",--14488
"111110001110001001110101100000000000",--14489
"001111010110000011000000000000000010",--14490
"111110010110001011000101100000000000",--14491
"111110010100000010110101000000000000",--14492
"001101010010000010110000000000000011",--14493
"011100010111000000000000000000000011",--14494
"101110010101111000000010100000000000",--14495
"011111010101000000110000000000010000",--14496
"000101000000000000000011100010110000",--14497
"111110001100001001110101100000000000",--14498
"001101010010000010110000000000001001",--14499
"001111010110000011000000000000000000",--14500
"111110010110001011000101100000000000",--14501
"111110010100000010110101000000000000",--14502
"111110001110001001010011100000000000",--14503
"001111010110000010110000000000000001",--14504
"111110001110001010110011100000000000",--14505
"111110010100000001110011100000000000",--14506
"111110001010001001100010100000000000",--14507
"001111010110000001100000000000000010",--14508
"111110001010001001100010100000000000",--14509
"111110001110000001010010100000000000",--14510
"011111010101000000110000000000000001",--14511
"111110001010010000010010100000000000",--14512
"111110010010001010010011000000000000",--14513
"111110010000001001010010100000000000",--14514
"111110001100010001010010100000000000",--14515
"010110001011000000000000000011110100",--14516
"001101010010000010010000000000000110",--14517
"011100010011000000000000000000000110",--14518
"111110001010100000000010100000000000",--14519
"111110010010010001010010100000000000",--14520
"001111010000000001100000000000000100",--14521
"111110001010001001100010100000000000",--14522
"001011000000000001010000000100101111",--14523
"000101000000000000000011100011000010",--14524
"111110001010100000000010100000000000",--14525
"111110010010000001010010100000000000",--14526
"001111010000000001100000000000000100",--14527
"111110001010001001100010100000000000",--14528
"001011000000000001010000000100101111",--14529
"001111000000000001010000000100101111",--14530
"101111001101110001101011110111001100",--14531
"101111001101100001101100110011001101",--14532
"010110001101000001010000000011100011",--14533
"001101001110000010000000000000000001",--14534
"010011010001000000000000000011100001",--14535
"001101010000000010000000000100110001",--14536
"001101010000000010010000000000000000",--14537
"010011010011000000000000000011001100",--14538
"001101010010000010100000000101101101",--14539
"001111000000000001010000000100101010",--14540
"001101010100000010110000000000000101",--14541
"001111010110000001100000000000000000",--14542
"111110001010010001100010100000000000",--14543
"001111000000000001100000000100101011",--14544
"001111010110000001110000000000000001",--14545
"111110001100010001110011000000000000",--14546
"001111000000000001110000000100101100",--14547
"001111010110000010000000000000000010",--14548
"111110001110010010000011100000000000",--14549
"001101010010000010110000000010111110",--14550
"001101010100000011000000000000000001",--14551
"011111011001000000010000000000111100",--14552
"001111010110000010000000000000000000",--14553
"111110010000010001010100000000000000",--14554
"001111010110000010010000000000000001",--14555
"111110010000001010010100000000000000",--14556
"001111000000000010010000000011111011",--14557
"111110010000001010010100100000000000",--14558
"111110010010000001100100100000000001",--14559
"001101010100000010100000000000000100",--14560
"001111010100000010100000000000000001",--14561
"010110010101000010010000000000000111",--14562
"001111000000000010010000000011111100",--14563
"111110010000001010010100100000000000",--14564
"111110010010000001110100100000000001",--14565
"001111010100000010100000000000000010",--14566
"010110010101000010010000000000000010",--14567
"001111010110000010010000000000000001",--14568
"011110010011000000000000000000101000",--14569
"001111010110000010000000000000000010",--14570
"111110010000010001100100000000000000",--14571
"001111010110000010010000000000000011",--14572
"111110010000001010010100000000000000",--14573
"001111000000000010010000000011111010",--14574
"111110010000001010010100100000000000",--14575
"111110010010000001010100100000000001",--14576
"001111010100000010100000000000000000",--14577
"010110010101000010010000000000000111",--14578
"001111000000000010010000000011111100",--14579
"111110010000001010010100100000000000",--14580
"111110010010000001110100100000000001",--14581
"001111010100000010100000000000000010",--14582
"010110010101000010010000000000000010",--14583
"001111010110000010010000000000000011",--14584
"011110010011000000000000000000010101",--14585
"001111010110000010000000000000000100",--14586
"111110010000010001110011100000000000",--14587
"001111010110000010000000000000000101",--14588
"111110001110001010000011100000000000",--14589
"001111000000000010000000000011111010",--14590
"111110001110001010000100000000000000",--14591
"111110010000000001010010100000000001",--14592
"001111010100000010000000000000000000",--14593
"010110010001000001010000000000000111",--14594
"001111000000000001010000000011111011",--14595
"111110001110001001010010100000000000",--14596
"111110001010000001100010100000000001",--14597
"001111010100000001100000000000000001",--14598
"010110001101000001010000000000000010",--14599
"001111010110000001010000000000000101",--14600
"011110001011000000000000000000000010",--14601
"101000000001111000000101000000000000",--14602
"000101000000000000000011100101100101",--14603
"001011000000000001110000000100101111",--14604
"101001000000000010100000000000000011",--14605
"000101000000000000000011100101100101",--14606
"001011000000000010000000000100101111",--14607
"101001000000000010100000000000000010",--14608
"000101000000000000000011100101100101",--14609
"001011000000000010000000000100101111",--14610
"101001000000000010100000000000000001",--14611
"000101000000000000000011100101100101",--14612
"011111011001000000100000000000001111",--14613
"001111010110000010000000000000000000",--14614
"011010010001000000000000000000001011",--14615
"001111010110000010000000000000000001",--14616
"111110010000001001010010100000000000",--14617
"001111010110000010000000000000000010",--14618
"111110010000001001100011000000000000",--14619
"111110001010000001100010100000000000",--14620
"001111010110000001100000000000000011",--14621
"111110001100001001110011000000000000",--14622
"111110001010000001100010100000000000",--14623
"001011000000000001010000000100101111",--14624
"101001000000000010100000000000000001",--14625
"000101000000000000000011100101100101",--14626
"101000000001111000000101000000000000",--14627
"000101000000000000000011100101100101",--14628
"001111010110000010000000000000000000",--14629
"011110010001000000000000000000000010",--14630
"101000000001111000000101000000000000",--14631
"000101000000000000000011100101100101",--14632
"001111010110000010010000000000000001",--14633
"111110010010001001010100100000000000",--14634
"001111010110000010100000000000000010",--14635
"111110010100001001100101000000000000",--14636
"111110010010000010100100100000000000",--14637
"001111010110000010100000000000000011",--14638
"111110010100001001110101000000000000",--14639
"111110010010000010100100100000000000",--14640
"111110001010001001010101000000000000",--14641
"001101010100000011010000000000000100",--14642
"001111011010000010110000000000000000",--14643
"111110010100001010110101000000000000",--14644
"111110001100001001100101100000000000",--14645
"001111011010000011000000000000000001",--14646
"111110010110001011000101100000000000",--14647
"111110010100000010110101000000000000",--14648
"111110001110001001110101100000000000",--14649
"001111011010000011000000000000000010",--14650
"111110010110001011000101100000000000",--14651
"111110010100000010110101000000000000",--14652
"001101010100000011010000000000000011",--14653
"011100011011000000000000000000000011",--14654
"101110010101111000000010100000000000",--14655
"011111011001000000110000000000010000",--14656
"000101000000000000000011100101010000",--14657
"111110001100001001110101100000000000",--14658
"001101010100000011010000000000001001",--14659
"001111011010000011000000000000000000",--14660
"111110010110001011000101100000000000",--14661
"111110010100000010110101000000000000",--14662
"111110001110001001010011100000000000",--14663
"001111011010000010110000000000000001",--14664
"111110001110001010110011100000000000",--14665
"111110010100000001110011100000000000",--14666
"111110001010001001100010100000000000",--14667
"001111011010000001100000000000000010",--14668
"111110001010001001100010100000000000",--14669
"111110001110000001010010100000000000",--14670
"011111011001000000110000000000000001",--14671
"111110001010010000010010100000000000",--14672
"111110010010001010010011000000000000",--14673
"111110010000001001010010100000000000",--14674
"111110001100010001010010100000000000",--14675
"010110001011000000000000000000001111",--14676
"001101010100000010100000000000000110",--14677
"011100010101000000000000000000000110",--14678
"111110001010100000000010100000000000",--14679
"111110010010010001010010100000000000",--14680
"001111010110000001100000000000000100",--14681
"111110001010001001100010100000000000",--14682
"001011000000000001010000000100101111",--14683
"000101000000000000000011100101100010",--14684
"111110001010100000000010100000000000",--14685
"111110010010000001010010100000000000",--14686
"001111010110000001100000000000000100",--14687
"111110001010001001100010100000000000",--14688
"001011000000000001010000000100101111",--14689
"101001000000000010100000000000000001",--14690
"000101000000000000000011100101100101",--14691
"101000000001111000000101000000000000",--14692
"001111000000000001010000000100101111",--14693
"010000010101000000000000000000100101",--14694
"101111001101110001101011111001001100",--14695
"101111001101100001101100110011001101",--14696
"010110001101000001010000000000100010",--14697
"101111001101110001100011110000100011",--14698
"101111001101100001101101011100001010",--14699
"111110001010000001100010100000000000",--14700
"001111000000000001100000000101100100",--14701
"111110001100001001010011000000000000",--14702
"001111000000000001110000000100101010",--14703
"111110001100000001110011000000000000",--14704
"001111000000000001110000000101100101",--14705
"111110001110001001010011100000000000",--14706
"001111000000000010000000000100101011",--14707
"111110001110000010000011100000000000",--14708
"001111000000000010000000000101100110",--14709
"111110010000001001010010100000000000",--14710
"001111000000000010000000000100101100",--14711
"111110001010000010000010100000000000",--14712
"001001111100000010001111111111110011",--14713
"101000010001111000000001000000000000",--14714
"101000000001111000000000100000000000",--14715
"101110001111111000000010000000000000",--14716
"101110001101111000000001100000000000",--14717
"001001111100000111111111111111110010",--14718
"101001111100010111100000000000001111",--14719
"000111000000000000000000011110001000",--14720
"101001111100000111100000000000001111",--14721
"001101111100000111111111111111110010",--14722
"011100000011000000000000000000101110",--14723
"101001000000000000010000000000000001",--14724
"001101111100000000101111111111110011",--14725
"101001111100010111100000000000001111",--14726
"000111000000000000000000100011100001",--14727
"101001111100000111100000000000001111",--14728
"001101111100000111111111111111110010",--14729
"011100000011000000000000000000100111",--14730
"000101000000000000000011100110010111",--14731
"001101010010000010010000000101101101",--14732
"001101010010000010010000000000000110",--14733
"010000010011000000000000000000001000",--14734
"101000010001111000000001000000000000",--14735
"101001000000000000010000000000000001",--14736
"001001111100000111111111111111110011",--14737
"101001111100010111100000000000001110",--14738
"000111000000000000000000100011100001",--14739
"101001111100000111100000000000001110",--14740
"001101111100000111111111111111110011",--14741
"011100000011000000000000000000011011",--14742
"001101111100000000011111111111110101",--14743
"001101000010000000100000000000000010",--14744
"010011000101000000000000000000001111",--14745
"001101000100000000100000000100110001",--14746
"101000000001111000000000100000000000",--14747
"001001111100000111111111111111110011",--14748
"101001111100010111100000000000001110",--14749
"000111000000000000000000100011100001",--14750
"101001111100000111100000000000001110",--14751
"001101111100000111111111111111110011",--14752
"011100000011000000000000000000010000",--14753
"101001000000000000010000000000000011",--14754
"001101111100000000101111111111110101",--14755
"101001111100010111100000000000001110",--14756
"000111000000000000000000110101111110",--14757
"101001111100000111100000000000001110",--14758
"001101111100000111111111111111110011",--14759
"011100000011000000000000000000001001",--14760
"101001000000000000010000000000000001",--14761
"001101111100000000101111111111110100",--14762
"001001111100000111111111111111110011",--14763
"101001111100010111100000000000001110",--14764
"000111000000000000000000111111111011",--14765
"101001111100000111100000000000001110",--14766
"001101111100000111111111111111110011",--14767
"011100000011000000000000000100100100",--14768
"000101000000000000000011101010011110",--14769
"001101111100000000011111111111110101",--14770
"001101000010000000100000000000000001",--14771
"010011000101000000000000000011100001",--14772
"001101000100000000100000000100110001",--14773
"001101000100000000110000000000000000",--14774
"010011000111000000000000000011001100",--14775
"001101000110000001000000000101101101",--14776
"001111000000000000110000000100101010",--14777
"001101001000000001010000000000000101",--14778
"001111001010000001000000000000000000",--14779
"111110000110010001000001100000000000",--14780
"001111000000000001000000000100101011",--14781
"001111001010000001010000000000000001",--14782
"111110001000010001010010000000000000",--14783
"001111000000000001010000000100101100",--14784
"001111001010000001100000000000000010",--14785
"111110001010010001100010100000000000",--14786
"001101000110000001010000000010111110",--14787
"001101001000000001100000000000000001",--14788
"011111001101000000010000000000111100",--14789
"001111001010000001100000000000000000",--14790
"111110001100010000110011000000000000",--14791
"001111001010000001110000000000000001",--14792
"111110001100001001110011000000000000",--14793
"001111000000000001110000000011111011",--14794
"111110001100001001110011100000000000",--14795
"111110001110000001000011100000000001",--14796
"001101001000000001000000000000000100",--14797
"001111001000000010000000000000000001",--14798
"010110010001000001110000000000000111",--14799
"001111000000000001110000000011111100",--14800
"111110001100001001110011100000000000",--14801
"111110001110000001010011100000000001",--14802
"001111001000000010000000000000000010",--14803
"010110010001000001110000000000000010",--14804
"001111001010000001110000000000000001",--14805
"011110001111000000000000000000101000",--14806
"001111001010000001100000000000000010",--14807
"111110001100010001000011000000000000",--14808
"001111001010000001110000000000000011",--14809
"111110001100001001110011000000000000",--14810
"001111000000000001110000000011111010",--14811
"111110001100001001110011100000000000",--14812
"111110001110000000110011100000000001",--14813
"001111001000000010000000000000000000",--14814
"010110010001000001110000000000000111",--14815
"001111000000000001110000000011111100",--14816
"111110001100001001110011100000000000",--14817
"111110001110000001010011100000000001",--14818
"001111001000000010000000000000000010",--14819
"010110010001000001110000000000000010",--14820
"001111001010000001110000000000000011",--14821
"011110001111000000000000000000010101",--14822
"001111001010000001100000000000000100",--14823
"111110001100010001010010100000000000",--14824
"001111001010000001100000000000000101",--14825
"111110001010001001100010100000000000",--14826
"001111000000000001100000000011111010",--14827
"111110001010001001100011000000000000",--14828
"111110001100000000110001100000000001",--14829
"001111001000000001100000000000000000",--14830
"010110001101000000110000000000000111",--14831
"001111000000000000110000000011111011",--14832
"111110001010001000110001100000000000",--14833
"111110000110000001000001100000000001",--14834
"001111001000000001000000000000000001",--14835
"010110001001000000110000000000000010",--14836
"001111001010000000110000000000000101",--14837
"011110000111000000000000000000000010",--14838
"101000000001111000000010000000000000",--14839
"000101000000000000000011101001010010",--14840
"001011000000000001010000000100101111",--14841
"101001000000000001000000000000000011",--14842
"000101000000000000000011101001010010",--14843
"001011000000000001100000000100101111",--14844
"101001000000000001000000000000000010",--14845
"000101000000000000000011101001010010",--14846
"001011000000000001100000000100101111",--14847
"101001000000000001000000000000000001",--14848
"000101000000000000000011101001010010",--14849
"011111001101000000100000000000001111",--14850
"001111001010000001100000000000000000",--14851
"011010001101000000000000000000001011",--14852
"001111001010000001100000000000000001",--14853
"111110001100001000110001100000000000",--14854
"001111001010000001100000000000000010",--14855
"111110001100001001000010000000000000",--14856
"111110000110000001000001100000000000",--14857
"001111001010000001000000000000000011",--14858
"111110001000001001010010000000000000",--14859
"111110000110000001000001100000000000",--14860
"001011000000000000110000000100101111",--14861
"101001000000000001000000000000000001",--14862
"000101000000000000000011101001010010",--14863
"101000000001111000000010000000000000",--14864
"000101000000000000000011101001010010",--14865
"001111001010000001100000000000000000",--14866
"011110001101000000000000000000000010",--14867
"101000000001111000000010000000000000",--14868
"000101000000000000000011101001010010",--14869
"001111001010000001110000000000000001",--14870
"111110001110001000110011100000000000",--14871
"001111001010000010000000000000000010",--14872
"111110010000001001000100000000000000",--14873
"111110001110000010000011100000000000",--14874
"001111001010000010000000000000000011",--14875
"111110010000001001010100000000000000",--14876
"111110001110000010000011100000000000",--14877
"111110000110001000110100000000000000",--14878
"001101001000000001110000000000000100",--14879
"001111001110000010010000000000000000",--14880
"111110010000001010010100000000000000",--14881
"111110001000001001000100100000000000",--14882
"001111001110000010100000000000000001",--14883
"111110010010001010100100100000000000",--14884
"111110010000000010010100000000000000",--14885
"111110001010001001010100100000000000",--14886
"001111001110000010100000000000000010",--14887
"111110010010001010100100100000000000",--14888
"111110010000000010010100000000000000",--14889
"001101001000000001110000000000000011",--14890
"011100001111000000000000000000000011",--14891
"101110010001111000000001100000000000",--14892
"011111001101000000110000000000010000",--14893
"000101000000000000000011101000111101",--14894
"111110001000001001010100100000000000",--14895
"001101001000000001110000000000001001",--14896
"001111001110000010100000000000000000",--14897
"111110010010001010100100100000000000",--14898
"111110010000000010010100000000000000",--14899
"111110001010001000110010100000000000",--14900
"001111001110000010010000000000000001",--14901
"111110001010001010010010100000000000",--14902
"111110010000000001010010100000000000",--14903
"111110000110001001000001100000000000",--14904
"001111001110000001000000000000000010",--14905
"111110000110001001000001100000000000",--14906
"111110001010000000110001100000000000",--14907
"011111001101000000110000000000000001",--14908
"111110000110010000010001100000000000",--14909
"111110001110001001110010000000000000",--14910
"111110001100001000110001100000000000",--14911
"111110001000010000110001100000000000",--14912
"010110000111000000000000000000001111",--14913
"001101001000000001000000000000000110",--14914
"011100001001000000000000000000000110",--14915
"111110000110100000000001100000000000",--14916
"111110001110010000110001100000000000",--14917
"001111001010000001000000000000000100",--14918
"111110000110001001000001100000000000",--14919
"001011000000000000110000000100101111",--14920
"000101000000000000000011101001001111",--14921
"111110000110100000000001100000000000",--14922
"111110001110000000110001100000000000",--14923
"001111001010000001000000000000000100",--14924
"111110000110001001000001100000000000",--14925
"001011000000000000110000000100101111",--14926
"101001000000000001000000000000000001",--14927
"000101000000000000000011101001010010",--14928
"101000000001111000000010000000000000",--14929
"001111000000000000110000000100101111",--14930
"010000001001000000000000000000100110",--14931
"101111001001110001001011111001001100",--14932
"101111001001100001001100110011001101",--14933
"010110001001000000110000000000100011",--14934
"101111001001110001000011110000100011",--14935
"101111001001100001001101011100001010",--14936
"111110000110000001000001100000000000",--14937
"001111000000000001000000000101100100",--14938
"111110001000001000110010000000000000",--14939
"001111000000000001010000000100101010",--14940
"111110001000000001010010000000000000",--14941
"001111000000000001010000000101100101",--14942
"111110001010001000110010100000000000",--14943
"001111000000000001100000000100101011",--14944
"111110001010000001100010100000000000",--14945
"001111000000000001100000000101100110",--14946
"111110001100001000110001100000000000",--14947
"001111000000000001100000000100101100",--14948
"111110000110000001100001100000000000",--14949
"001001111100000000101111111111110011",--14950
"101000000001111000000000100000000000",--14951
"101110001011111000001111100000000000",--14952
"101110000111111000000010100000000000",--14953
"101110001001111000000001100000000000",--14954
"101110111111111000000010000000000000",--14955
"001001111100000111111111111111110010",--14956
"101001111100010111100000000000001111",--14957
"000111000000000000000000011110001000",--14958
"101001111100000111100000000000001111",--14959
"001101111100000111111111111111110010",--14960
"011100000011000000000000000001100011",--14961
"101001000000000000010000000000000001",--14962
"001101111100000000101111111111110011",--14963
"101001111100010111100000000000001111",--14964
"000111000000000000000000100011100001",--14965
"101001111100000111100000000000001111",--14966
"001101111100000111111111111111110010",--14967
"011100000011000000000000000001011100",--14968
"000101000000000000000011101010000100",--14969
"001101000110000000110000000101101101",--14970
"001101000110000000110000000000000110",--14971
"010000000111000000000000000000000111",--14972
"101001000000000000010000000000000001",--14973
"001001111100000111111111111111110011",--14974
"101001111100010111100000000000001110",--14975
"000111000000000000000000100011100001",--14976
"101001111100000111100000000000001110",--14977
"001101111100000111111111111111110011",--14978
"011100000011000000000000000001010001",--14979
"001101111100000000011111111111110101",--14980
"001101000010000000100000000000000010",--14981
"010011000101000000000000000000001111",--14982
"001101000100000000100000000100110001",--14983
"101000000001111000000000100000000000",--14984
"001001111100000111111111111111110011",--14985
"101001111100010111100000000000001110",--14986
"000111000000000000000000100011100001",--14987
"101001111100000111100000000000001110",--14988
"001101111100000111111111111111110011",--14989
"011100000011000000000000000001000110",--14990
"101001000000000000010000000000000011",--14991
"001101111100000000101111111111110101",--14992
"101001111100010111100000000000001110",--14993
"000111000000000000000000110101111110",--14994
"101001111100000111100000000000001110",--14995
"001101111100000111111111111111110011",--14996
"011100000011000000000000000000111111",--14997
"101001000000000000010000000000000001",--14998
"001101111100000000101111111111110100",--14999
"001001111100000111111111111111110011",--15000
"101001111100010111100000000000001110",--15001
"000111000000000000000000111111111011",--15002
"101001111100000111100000000000001110",--15003
"001101111100000111111111111111110011",--15004
"011100000011000000000000000000110111",--15005
"001111000000000000110000000100100110",--15006
"001111000000000001000000000101100100",--15007
"111110000110001001000001100000000000",--15008
"001111000000000001000000000100100111",--15009
"001111000000000001010000000101100101",--15010
"111110001000001001010010000000000000",--15011
"111110000110000001000001100000000000",--15012
"001111000000000001000000000100101000",--15013
"001111000000000001010000000101100110",--15014
"111110001000001001010010000000000000",--15015
"111110000110000001000001100000000010",--15016
"001111111100000001001111111111111001",--15017
"111110000110001001000001100000000000",--15018
"001101111100000000101111111111111101",--15019
"001111000100000001010000000000000000",--15020
"001111000000000001100000000101100100",--15021
"111110001010001001100010100000000000",--15022
"001111000100000001100000000000000001",--15023
"001111000000000001110000000101100101",--15024
"111110001100001001110011000000000000",--15025
"111110001010000001100010100000000000",--15026
"001111000100000001100000000000000010",--15027
"001111000000000001110000000101100110",--15028
"111110001100001001110011000000000000",--15029
"111110001010000001100010100000000010",--15030
"010110000111000000000000000000001111",--15031
"001111000000000001100000000100011101",--15032
"001111000000000001110000000100100011",--15033
"111110000110001001110011100000000000",--15034
"111110001100000001110011000000000000",--15035
"001011000000000001100000000100011101",--15036
"001111000000000001100000000100011110",--15037
"001111000000000001110000000100100100",--15038
"111110000110001001110011100000000000",--15039
"111110001100000001110011000000000000",--15040
"001011000000000001100000000100011110",--15041
"001111000000000001100000000100011111",--15042
"001111000000000001110000000100100101",--15043
"111110000110001001110001100000000000",--15044
"111110001100000000110001100000000000",--15045
"001011000000000000110000000100011111",--15046
"010110001011000000000000000000001101",--15047
"111110001010001001010001100000000000",--15048
"111110000110001000110001100000000000",--15049
"001111111100000001011111111111110110",--15050
"111110000110001001010001100000000000",--15051
"001111000000000001100000000100011101",--15052
"111110001100000000110011000000000000",--15053
"001011000000000001100000000100011101",--15054
"001111000000000001100000000100011110",--15055
"111110001100000000110011000000000000",--15056
"001011000000000001100000000100011110",--15057
"001111000000000001100000000100011111",--15058
"111110001100000000110001100000000000",--15059
"001011000000000000110000000100011111",--15060
"001111000000000000110000000100101010",--15061
"001011000000000000110000000100010010",--15062
"001111000000000000110000000100101011",--15063
"001011000000000000110000000100010011",--15064
"001111000000000000110000000100101100",--15065
"001011000000000000110000000100010100",--15066
"001101000000000000010000000110101010",--15067
"101001000010010000010000000000000001",--15068
"010111000011000000000000000010010001",--15069
"001101000010000000100000000101101101",--15070
"001101000100000000110000000000001010",--15071
"001101000100000001000000000000000001",--15072
"001111000000000000110000000100101010",--15073
"001101000100000001010000000000000101",--15074
"001111001010000001000000000000000000",--15075
"111110000110010001000001100000000000",--15076
"001011000110000000110000000000000000",--15077
"001111000000000000110000000100101011",--15078
"001111001010000001000000000000000001",--15079
"111110000110010001000001100000000000",--15080
"001011000110000000110000000000000001",--15081
"001111000000000000110000000100101100",--15082
"001111001010000001000000000000000010",--15083
"111110000110010001000001100000000000",--15084
"001011000110000000110000000000000010",--15085
"011111001001000000100000000000001110",--15086
"001101000100000000100000000000000100",--15087
"001111000110000000110000000000000000",--15088
"001111000110000001000000000000000001",--15089
"001111000110000001010000000000000010",--15090
"001111000100000001100000000000000000",--15091
"111110001100001000110001100000000000",--15092
"001111000100000001100000000000000001",--15093
"111110001100001001000010000000000000",--15094
"111110000110000001000001100000000000",--15095
"001111000100000001000000000000000010",--15096
"111110001000001001010010000000000000",--15097
"111110000110000001000001100000000000",--15098
"001011000110000000110000000000000011",--15099
"000101000000000000000011101100100010",--15100
"010111001001000000100000000000100100",--15101
"001111000110000000110000000000000000",--15102
"001111000110000001000000000000000001",--15103
"001111000110000001010000000000000010",--15104
"111110000110001000110011000000000000",--15105
"001101000100000001010000000000000100",--15106
"001111001010000001110000000000000000",--15107
"111110001100001001110011000000000000",--15108
"111110001000001001000011100000000000",--15109
"001111001010000010000000000000000001",--15110
"111110001110001010000011100000000000",--15111
"111110001100000001110011000000000000",--15112
"111110001010001001010011100000000000",--15113
"001111001010000010000000000000000010",--15114
"111110001110001010000011100000000000",--15115
"111110001100000001110011000000000000",--15116
"001101000100000001010000000000000011",--15117
"011100001011000000000000000000000011",--15118
"101110001101111000000001100000000000",--15119
"011111001001000000110000000000010000",--15120
"000101000000000000000011101100100000",--15121
"111110001000001001010011100000000000",--15122
"001101000100000000100000000000001001",--15123
"001111000100000010000000000000000000",--15124
"111110001110001010000011100000000000",--15125
"111110001100000001110011000000000000",--15126
"111110001010001000110010100000000000",--15127
"001111000100000001110000000000000001",--15128
"111110001010001001110010100000000000",--15129
"111110001100000001010010100000000000",--15130
"111110000110001001000001100000000000",--15131
"001111000100000001000000000000000010",--15132
"111110000110001001000001100000000000",--15133
"111110001010000000110001100000000000",--15134
"011111001001000000110000000000000001",--15135
"111110000110010000010001100000000000",--15136
"001011000110000000110000000000000011",--15137
"101001000010010000010000000000000001",--15138
"010111000011000000000000000001001011",--15139
"001101000010000000100000000101101101",--15140
"001101000100000000110000000000001010",--15141
"001101000100000001000000000000000001",--15142
"001111000000000000110000000100101010",--15143
"001101000100000001010000000000000101",--15144
"001111001010000001000000000000000000",--15145
"111110000110010001000001100000000000",--15146
"001011000110000000110000000000000000",--15147
"001111000000000000110000000100101011",--15148
"001111001010000001000000000000000001",--15149
"111110000110010001000001100000000000",--15150
"001011000110000000110000000000000001",--15151
"001111000000000000110000000100101100",--15152
"001111001010000001000000000000000010",--15153
"111110000110010001000001100000000000",--15154
"001011000110000000110000000000000010",--15155
"011111001001000000100000000000001110",--15156
"001101000100000000100000000000000100",--15157
"001111000110000000110000000000000000",--15158
"001111000110000001000000000000000001",--15159
"001111000110000001010000000000000010",--15160
"001111000100000001100000000000000000",--15161
"111110001100001000110001100000000000",--15162
"001111000100000001100000000000000001",--15163
"111110001100001001000010000000000000",--15164
"111110000110000001000001100000000000",--15165
"001111000100000001000000000000000010",--15166
"111110001000001001010010000000000000",--15167
"111110000110000001000001100000000000",--15168
"001011000110000000110000000000000011",--15169
"000101000000000000000011101101101000",--15170
"010111001001000000100000000000100100",--15171
"001111000110000000110000000000000000",--15172
"001111000110000001000000000000000001",--15173
"001111000110000001010000000000000010",--15174
"111110000110001000110011000000000000",--15175
"001101000100000001010000000000000100",--15176
"001111001010000001110000000000000000",--15177
"111110001100001001110011000000000000",--15178
"111110001000001001000011100000000000",--15179
"001111001010000010000000000000000001",--15180
"111110001110001010000011100000000000",--15181
"111110001100000001110011000000000000",--15182
"111110001010001001010011100000000000",--15183
"001111001010000010000000000000000010",--15184
"111110001110001010000011100000000000",--15185
"111110001100000001110011000000000000",--15186
"001101000100000001010000000000000011",--15187
"011100001011000000000000000000000011",--15188
"101110001101111000000001100000000000",--15189
"011111001001000000110000000000010000",--15190
"000101000000000000000011101101100110",--15191
"111110001000001001010011100000000000",--15192
"001101000100000000100000000000001001",--15193
"001111000100000010000000000000000000",--15194
"111110001110001010000011100000000000",--15195
"111110001100000001110011000000000000",--15196
"111110001010001000110010100000000000",--15197
"001111000100000001110000000000000001",--15198
"111110001010001001110010100000000000",--15199
"111110001100000001010010100000000000",--15200
"111110000110001001000001100000000000",--15201
"001111000100000001000000000000000010",--15202
"111110000110001001000001100000000000",--15203
"111110001010000000110001100000000000",--15204
"011111001001000000110000000000000001",--15205
"111110000110010000010001100000000000",--15206
"001011000110000000110000000000000011",--15207
"101001000010010000100000000000000001",--15208
"101001000000000000010000000100101010",--15209
"001001111100000111111111111111110101",--15210
"101001111100010111100000000000001100",--15211
"000111000000000000000000011001101110",--15212
"101001111100000111100000000000001100",--15213
"001101111100000111111111111111110101",--15214
"001101000000000000010000000000000011",--15215
"101001000010010000010000000000000001",--15216
"010111000011000000000000000011101001",--15217
"001101000010000000100000000000000100",--15218
"001101000100000000110000000000000001",--15219
"101111000111110000110100111001101110",--15220
"101111000111100000110110101100101000",--15221
"001011000000000000110000000100101101",--15222
"001101000000000001000000000100110000",--15223
"001101001000000001010000000000000000",--15224
"001101001010000001100000000000000000",--15225
"001001111100000000011111111111110101",--15226
"001001111100000000111111111111110100",--15227
"001001111100000000101111111111110011",--15228
"010011001101000000000000000010000000",--15229
"001001111100000001001111111111110010",--15230
"011111001101011000110000000000001000",--15231
"101000001011111000000001000000000000",--15232
"101001000000000000010000000000000001",--15233
"001001111100000111111111111111110001",--15234
"101001111100010111100000000000010000",--15235
"000111000000000000000010101111001101",--15236
"101001111100000111100000000000010000",--15237
"001101111100000111111111111111110001",--15238
"000101000000000000000011101111110110",--15239
"001101001100000001110000000101101101",--15240
"001101001110000010000000000000001010",--15241
"001111010000000000110000000000000000",--15242
"001111010000000001000000000000000001",--15243
"001111010000000001010000000000000010",--15244
"001101000110000010010000000000000001",--15245
"001100010010000001100011000000000000",--15246
"001101001110000010010000000000000001",--15247
"011111010011000000010000000000111000",--15248
"001101000110000010000000000000000000",--15249
"001111001100000001100000000000000000",--15250
"111110001100010000110011000000000000",--15251
"001111001100000001110000000000000001",--15252
"111110001100001001110011000000000000",--15253
"001111010000000001110000000000000001",--15254
"111110001100001001110011100000000000",--15255
"111110001110000001000011100000000001",--15256
"001101001110000001110000000000000100",--15257
"001111001110000010000000000000000001",--15258
"010110010001000001110000000000000111",--15259
"001111010000000001110000000000000010",--15260
"111110001100001001110011100000000000",--15261
"111110001110000001010011100000000001",--15262
"001111001110000010000000000000000010",--15263
"010110010001000001110000000000000010",--15264
"001111001100000001110000000000000001",--15265
"011110001111000000000000000000100100",--15266
"001111001100000001100000000000000010",--15267
"111110001100010001000011000000000000",--15268
"001111001100000001110000000000000011",--15269
"111110001100001001110011000000000000",--15270
"001111010000000001110000000000000000",--15271
"111110001100001001110011100000000000",--15272
"111110001110000000110011100000000001",--15273
"001111001110000010000000000000000000",--15274
"010110010001000001110000000000000111",--15275
"001111010000000001110000000000000010",--15276
"111110001100001001110011100000000000",--15277
"111110001110000001010011100000000001",--15278
"001111001110000010000000000000000010",--15279
"010110010001000001110000000000000010",--15280
"001111001100000001110000000000000011",--15281
"011110001111000000000000000000010010",--15282
"001111001100000001100000000000000100",--15283
"111110001100010001010010100000000000",--15284
"001111001100000001100000000000000101",--15285
"111110001010001001100010100000000000",--15286
"001111010000000001100000000000000000",--15287
"111110001010001001100011000000000000",--15288
"111110001100000000110001100000000001",--15289
"001111001110000001100000000000000000",--15290
"010110001101000000110000000000111010",--15291
"001111010000000000110000000000000001",--15292
"111110001010001000110001100000000000",--15293
"111110000110000001000001100000000001",--15294
"001111001110000001000000000000000001",--15295
"010110001001000000110000000000110101",--15296
"001111001100000000110000000000000101",--15297
"010010000111000000000000000000110011",--15298
"001011000000000001010000000100101111",--15299
"000101000000000000000011101111101100",--15300
"001011000000000001100000000100101111",--15301
"000101000000000000000011101111101100",--15302
"001011000000000001100000000100101111",--15303
"000101000000000000000011101111101100",--15304
"011111010011000000100000000000000110",--15305
"001111001100000000110000000000000000",--15306
"011010000111000000000000000000101010",--15307
"001111010000000001000000000000000011",--15308
"111110000110001001000001100000000000",--15309
"001011000000000000110000000100101111",--15310
"000101000000000000000011101111101100",--15311
"001111001100000001100000000000000000",--15312
"010010001101000000000000000000100100",--15313
"001111001100000001110000000000000001",--15314
"111110001110001000110001100000000000",--15315
"001111001100000001110000000000000010",--15316
"111110001110001001000010000000000000",--15317
"111110000110000001000001100000000000",--15318
"001111001100000001000000000000000011",--15319
"111110001000001001010010000000000000",--15320
"111110000110000001000001100000000000",--15321
"001111010000000001000000000000000011",--15322
"111110000110001000110010100000000000",--15323
"111110001100001001000010000000000000",--15324
"111110001010010001000010000000000000",--15325
"010110001001000000000000000000010111",--15326
"001101001110000001110000000000000110",--15327
"011100001111000000000000000000000110",--15328
"111110001000100000000010000000000000",--15329
"111110000110010001000001100000000000",--15330
"001111001100000001000000000000000100",--15331
"111110000110001001000001100000000000",--15332
"001011000000000000110000000100101111",--15333
"000101000000000000000011101111101100",--15334
"111110001000100000000010000000000000",--15335
"111110000110000001000001100000000000",--15336
"001111001100000001000000000000000100",--15337
"111110000110001001000001100000000000",--15338
"001011000000000000110000000100101111",--15339
"001111000000000000110000000100101111",--15340
"001111000000000001000000000100101101",--15341
"010110001001000000110000000000000111",--15342
"101000001011111000000001000000000000",--15343
"101001000000000000010000000000000001",--15344
"001001111100000111111111111111110001",--15345
"101001111100010111100000000000010000",--15346
"000111000000000000000010101111001101",--15347
"101001111100000111100000000000010000",--15348
"001101111100000111111111111111110001",--15349
"101001000000000000010000000000000001",--15350
"001101111100000000101111111111110010",--15351
"001101111100000000111111111111110100",--15352
"001001111100000111111111111111110001",--15353
"101001111100010111100000000000010000",--15354
"000111000000000000000010110111111111",--15355
"101001111100000111100000000000010000",--15356
"001101111100000111111111111111110001",--15357
"001111000000000000110000000100101101",--15358
"101111001001110001001011110111001100",--15359
"101111001001100001001100110011001101",--15360
"010110000111000001000000000001001111",--15361
"101111001001110001000100110010111110",--15362
"101111001001100001001011110000100000",--15363
"010110001001000000110000000001001100",--15364
"001101000000000000010000000100101001",--15365
"101000000011000000010000100010000010",--15366
"001101000000000000100000000100101110",--15367
"101000000010000000100000100000000000",--15368
"001101111100000000101111111111110011",--15369
"001101000100000000110000000000000000",--15370
"011100000011000000110000000001000101",--15371
"101000000001111000000000100000000000",--15372
"001101000000000000100000000100110000",--15373
"001001111100000111111111111111110010",--15374
"101001111100010111100000000000001111",--15375
"000111000000000000000000111111111011",--15376
"101001111100000111100000000000001111",--15377
"001101111100000111111111111111110010",--15378
"011100000011000000000000000000111101",--15379
"001101111100000000011111111111110100",--15380
"001101000010000000010000000000000000",--15381
"001111000000000000110000000100100110",--15382
"001111000010000001000000000000000000",--15383
"111110000110001001000001100000000000",--15384
"001111000000000001000000000100100111",--15385
"001111000010000001010000000000000001",--15386
"111110001000001001010010000000000000",--15387
"111110000110000001000001100000000000",--15388
"001111000000000001000000000100101000",--15389
"001111000010000001010000000000000010",--15390
"111110001000001001010010000000000000",--15391
"111110000110000001000001100000000000",--15392
"001101111100000000101111111111110011",--15393
"001111000100000001000000000000000010",--15394
"001111111100000001011111111111111001",--15395
"111110001000001001010011000000000000",--15396
"111110001100001000110001100000000000",--15397
"001101111100000000101111111111111101",--15398
"001111000100000001100000000000000000",--15399
"001111000010000001110000000000000000",--15400
"111110001100001001110011000000000000",--15401
"001111000100000001110000000000000001",--15402
"001111000010000010000000000000000001",--15403
"111110001110001010000011100000000000",--15404
"111110001100000001110011000000000000",--15405
"001111000100000001110000000000000010",--15406
"001111000010000010000000000000000010",--15407
"111110001110001010000011100000000000",--15408
"111110001100000001110011000000000000",--15409
"111110001000001001100010000000000000",--15410
"010110000111000000000000000000001111",--15411
"001111000000000001100000000100011101",--15412
"001111000000000001110000000100100011",--15413
"111110000110001001110011100000000000",--15414
"111110001100000001110011000000000000",--15415
"001011000000000001100000000100011101",--15416
"001111000000000001100000000100011110",--15417
"001111000000000001110000000100100100",--15418
"111110000110001001110011100000000000",--15419
"111110001100000001110011000000000000",--15420
"001011000000000001100000000100011110",--15421
"001111000000000001100000000100011111",--15422
"001111000000000001110000000100100101",--15423
"111110000110001001110001100000000000",--15424
"111110001100000000110001100000000000",--15425
"001011000000000000110000000100011111",--15426
"010110001001000000000000000000001101",--15427
"111110001000001001000001100000000000",--15428
"111110000110001000110001100000000000",--15429
"001111111100000001001111111111110110",--15430
"111110000110001001000001100000000000",--15431
"001111000000000001100000000100011101",--15432
"111110001100000000110011000000000000",--15433
"001011000000000001100000000100011101",--15434
"001111000000000001100000000100011110",--15435
"111110001100000000110011000000000000",--15436
"001011000000000001100000000100011110",--15437
"001111000000000001100000000100011111",--15438
"111110001100000000110001100000000000",--15439
"001011000000000000110000000100011111",--15440
"001101111100000000011111111111110101",--15441
"101001000010010000010000000000000001",--15442
"001111111100000000111111111111111001",--15443
"001111111100000001001111111111110110",--15444
"001101111100000000101111111111111101",--15445
"001001111100000111111111111111110010",--15446
"101001111100010111100000000000001111",--15447
"000111000000000000000011001000010100",--15448
"101001111100000111100000000000001111",--15449
"001101111100000111111111111111110010",--15450
"101111000111110000110011110111001100",--15451
"101111000111100000111100110011001101",--15452
"001111111100000001001111111111111110",--15453
"010110001000000000111111100000000000",--15454
"001101111100000000011111111111111010",--15455
"001101000010000000010000000000000010",--15456
"001101111100000000101111111111111011",--15457
"011011000101000001000000000000000100",--15458
"101001000100000000110000000000000001",--15459
"101001000000000001001111111111111111",--15460
"001101111100000001011111111111111100",--15461
"001000001010000000110010000000000000",--15462
"011111000010000000101111100000000000",--15463
"001101111100000000011111111111111000",--15464
"001111000010000000110000000000000000",--15465
"111110000110010000010001100000000010",--15466
"111110001000001000110001100000000000",--15467
"101001000100000000010000000000000001",--15468
"001111000000000001000000000100101101",--15469
"001111111100000001010000000000000000",--15470
"111110001010000001000010000000000000",--15471
"001101111100000000101111111111111101",--15472
"001101111100000000111111111111111111",--15473
"011011000010000001011111100000000000",--15474
"000101000000000000000011010111010000",--15475
"101111001001110001000100111001101110",--15476
"101111001001100001000110101100101000",--15477
"001011000000000001000000000100101101",--15478
"001101000000000000100000000100110000",--15479
"001011111100000000110000000000000000",--15480
"001001111100000000011111111111111111",--15481
"101000000011111000000001100000000000",--15482
"101000000001111000000000100000000000",--15483
"001001111100000111111111111111111110",--15484
"101001111100010111100000000000000011",--15485
"000111000000000000000010110111111111",--15486
"101001111100000111100000000000000011",--15487
"001101111100000111111111111111111110",--15488
"001111000000000000110000000100101101",--15489
"101111001001110001001011110111001100",--15490
"101111001001100001001100110011001101",--15491
"010110000110000001001111100000000000",--15492
"101111001001110001000100110010111110",--15493
"101111001001100001001011110000100000",--15494
"010110001000000000111111100000000000",--15495
"001101000000000000010000000100101001",--15496
"001101000010000000010000000101101101",--15497
"001101000010000000100000000000000001",--15498
"011111000101000000010000000000010011",--15499
"001101111100000000101111111111111111",--15500
"001101000100000000100000000000000000",--15501
"001101000000000000110000000100101110",--15502
"001011000000000000000000000100100110",--15503
"001011000000000000000000000100100111",--15504
"001011000000000000000000000100101000",--15505
"101001000110010001000000000000000001",--15506
"101001000110010000110000000000000001",--15507
"001110000100000000110001100000000000",--15508
"011110000111000000000000000000000010",--15509
"101110000001111000000001100000000000",--15510
"000101000000000000000011110010011100",--15511
"010110000111000000000000000000000010",--15512
"101110000011111000000001100000000000",--15513
"000101000000000000000011110010011100",--15514
"101110000101111000000001100000000000",--15515
"101110000111111000000001100000000010",--15516
"001011001000000000110000000100100110",--15517
"000101000000000000000011110011110101",--15518
"011111000101000000100000000000001000",--15519
"001101000010000000100000000000000100",--15520
"001111000100010000110000000000000000",--15521
"001011000000000000110000000100100110",--15522
"001111000100010000110000000000000001",--15523
"001011000000000000110000000100100111",--15524
"001111000100010000110000000000000010",--15525
"001011000000000000110000000100101000",--15526
"000101000000000000000011110011110101",--15527
"001111000000000000110000000100101010",--15528
"001101000010000000100000000000000101",--15529
"001111000100000001000000000000000000",--15530
"111110000110010001000001100000000000",--15531
"001111000000000001000000000100101011",--15532
"001111000100000001010000000000000001",--15533
"111110001000010001010010000000000000",--15534
"001111000000000001010000000100101100",--15535
"001111000100000001100000000000000010",--15536
"111110001010010001100010100000000000",--15537
"001101000010000000100000000000000100",--15538
"001111000100000001100000000000000000",--15539
"111110000110001001100011000000000000",--15540
"001111000100000001110000000000000001",--15541
"111110001000001001110011100000000000",--15542
"001111000100000010000000000000000010",--15543
"111110001010001010000100000000000000",--15544
"001101000010000000100000000000000011",--15545
"011100000101000000000000000000000100",--15546
"001011000000000001100000000100100110",--15547
"001011000000000001110000000100100111",--15548
"001011000000000010000000000100101000",--15549
"000101000000000000000011110011011011",--15550
"001101000010000000100000000000001001",--15551
"001111000100000010010000000000000010",--15552
"111110001000001010010100100000000000",--15553
"001111000100000010100000000000000001",--15554
"111110001010001010100101000000000000",--15555
"111110010010000010100100100000000000",--15556
"101111000001110010100011111100000000",--15557
"111110010010001010100100100000000000",--15558
"111110001100000010010011000000000000",--15559
"001011000000000001100000000100100110",--15560
"001111000100000001100000000000000010",--15561
"111110000110001001100011000000000000",--15562
"001111000100000010010000000000000000",--15563
"111110001010001010010010100000000000",--15564
"111110001100000001010010100000000000",--15565
"101111000001110001100011111100000000",--15566
"111110001010001001100010100000000000",--15567
"111110001110000001010010100000000000",--15568
"001011000000000001010000000100100111",--15569
"001111000100000001010000000000000001",--15570
"111110000110001001010001100000000000",--15571
"001111000100000001010000000000000000",--15572
"111110001000001001010010000000000000",--15573
"111110000110000001000001100000000000",--15574
"101111000001110001000011111100000000",--15575
"111110000110001001000001100000000000",--15576
"111110010000000000110001100000000000",--15577
"001011000000000000110000000100101000",--15578
"001111000000000000110000000100100110",--15579
"111110000110001000110001100000000000",--15580
"001111000000000001000000000100100111",--15581
"111110001000001001000010000000000000",--15582
"111110000110000001000001100000000000",--15583
"001111000000000001000000000100101000",--15584
"111110001000001001000010000000000000",--15585
"111110000110000001000001100000000000",--15586
"111110000110100000000001100000000000",--15587
"011110000111000000000000000000000010",--15588
"101110000011111000000001100000000000",--15589
"000101000000000000000011110011101100",--15590
"001101000010000000100000000000000110",--15591
"011100000101000000000000000000000010",--15592
"111110000110011000000001100000000000",--15593
"000101000000000000000011110011101100",--15594
"111110000110011000000001100000000010",--15595
"001111000000000001000000000100100110",--15596
"111110001000001000110010000000000000",--15597
"001011000000000001000000000100100110",--15598
"001111000000000001000000000100100111",--15599
"111110001000001000110010000000000000",--15600
"001011000000000001000000000100100111",--15601
"001111000000000001000000000100101000",--15602
"111110001000001000110001100000000000",--15603
"001011000000000000110000000100101000",--15604
"001101000010000000100000000000000000",--15605
"001101000010000000110000000000001000",--15606
"001111000110000000110000000000000000",--15607
"001011000000000000110000000100100011",--15608
"001111000110000000110000000000000001",--15609
"001011000000000000110000000100100100",--15610
"001111000110000000110000000000000010",--15611
"001011000000000000110000000100100101",--15612
"001001111100000000011111111111111110",--15613
"011111000101000000010000000000100011",--15614
"001111000000000000110000000100101010",--15615
"001101000010000000100000000000000101",--15616
"001111000100000001000000000000000000",--15617
"111110000110010001000001100000000000",--15618
"101111001001110001000011110101001100",--15619
"101111001001100001001100110011001101",--15620
"111110000110001001000010000000000000",--15621
"101110001000110000000010000000000000",--15622
"101111000001110001010100000110100000",--15623
"111110001000001001010010000000000000",--15624
"111110000110010001000001100000000000",--15625
"101111000001110001000100000100100000",--15626
"001111000000000001010000000100101100",--15627
"001111000100000001100000000000000010",--15628
"111110001010010001100010100000000000",--15629
"101111001101110001100011110101001100",--15630
"101111001101100001101100110011001101",--15631
"111110001010001001100011000000000000",--15632
"101110001100110000000011000000000000",--15633
"101111000001110001110100000110100000",--15634
"111110001100001001110011000000000000",--15635
"111110001010010001100010100000000000",--15636
"101111000001110001100100000100100000",--15637
"010110001001000000110000000000000101",--15638
"010110001101000001010000000000000010",--15639
"101111000001110000110100001101111111",--15640
"000101000000000000000011110100100000",--15641
"101110000001111000000001100000000000",--15642
"000101000000000000000011110100100000",--15643
"010110001101000001010000000000000010",--15644
"101110000001111000000001100000000000",--15645
"000101000000000000000011110100100000",--15646
"101111000001110000110100001101111111",--15647
"001011000000000000110000000100100100",--15648
"000101000000000000000011111001000100",--15649
"011111000101000000100000000000001111",--15650
"001111000000000000110000000100101011",--15651
"101111000001110001000011111010000000",--15652
"111110000110001001000001100000000000",--15653
"001001111100000111111111111111111101",--15654
"000111000000000000000111011000000010",--15655
"001101111100000111111111111111111101",--15656
"111110000110001000110001100000000000",--15657
"101111000001110001000100001101111111",--15658
"111110001000001000110010000000000000",--15659
"001011000000000001000000000100100011",--15660
"101111000001110001000100001101111111",--15661
"111110000110010000010001100000000010",--15662
"111110001000001000110001100000000000",--15663
"001011000000000000110000000100100100",--15664
"000101000000000000000011111001000100",--15665
"011111000101000000110000000000011111",--15666
"001111000000000000110000000100101010",--15667
"001101000010000000100000000000000101",--15668
"001111000100000001000000000000000000",--15669
"111110000110010001000001100000000000",--15670
"001111000000000001000000000100101100",--15671
"001111000100000001010000000000000010",--15672
"111110001000010001010010000000000000",--15673
"111110000110001000110001100000000000",--15674
"111110001000001001000010000000000000",--15675
"111110000110000001000001100000000000",--15676
"111110000110100000000001100000000000",--15677
"101111001001110001000011110111001100",--15678
"101111001001100001001100110011001100",--15679
"111110000110001001000001100000000000",--15680
"101110000110110000000010000000000000",--15681
"111110000110010001000001100000000000",--15682
"101111001001110001000100000001001001",--15683
"101111001001100001000000111111011011",--15684
"111110000110001001000001100000000000",--15685
"001001111100000111111111111111111101",--15686
"000111000000000000000111010110111000",--15687
"001101111100000111111111111111111101",--15688
"111110000110001000110001100000000000",--15689
"101111000001110001000100001101111111",--15690
"111110000110001001000010000000000000",--15691
"001011000000000001000000000100100100",--15692
"111110000110010000010001100000000010",--15693
"101111000001110001000100001101111111",--15694
"111110000110001001000001100000000000",--15695
"001011000000000000110000000100100101",--15696
"000101000000000000000011111001000100",--15697
"011111000101000001000000000011110001",--15698
"001111000000000000110000000100101010",--15699
"001101000010000000100000000000000101",--15700
"001111000100000001000000000000000000",--15701
"111110000110010001000001100000000000",--15702
"001101000010000000110000000000000100",--15703
"001111000110000001000000000000000000",--15704
"111110001000100000000010000000000000",--15705
"111110000110001001000001100000000000",--15706
"001111000000000001000000000100101100",--15707
"001111000100000001010000000000000010",--15708
"111110001000010001010010000000000000",--15709
"001111000110000001010000000000000010",--15710
"111110001010100000000010100000000000",--15711
"111110001000001001010010000000000000",--15712
"111110000110001000110010100000000000",--15713
"111110001000001001000011000000000000",--15714
"111110001010000001100010100000000000",--15715
"101110000111111000000011000000000001",--15716
"101111001111110001110011100011010001",--15717
"101111001111100001111011011100010111",--15718
"010110001111000001100000000000000010",--15719
"101111000001110000110100000101110000",--15720
"000101000000000000000011110111000110",--15721
"111110000110011000000001100000000000",--15722
"111110001000001000110001100000000001",--15723
"010110000111000000010000000000000010",--15724
"101001000000000001000000000000000001",--15725
"000101000000000000000011110101110100",--15726
"011010000111000000100000000000000010",--15727
"101001000000000001001111111111111111",--15728
"000101000000000000000011110101110100",--15729
"101000000001111000000010000000000000",--15730
"000101000000000000000011110101110101",--15731
"111110000110011000000001100000000000",--15732
"111110000110001000110010000000000000",--15733
"101111000001110001100100001011110010",--15734
"111110001100001001000011000000000000",--15735
"101111001111110001110011110100110010",--15736
"101111001111100001110001011001000011",--15737
"111110001100001001110011000000000000",--15738
"101111000001110001110100001011001000",--15739
"111110001110001001000011100000000000",--15740
"101111000001110010000100000110101000",--15741
"111110010000000001100011000000000000",--15742
"111110001100011000000011000000000000",--15743
"111110001110001001100011000000000000",--15744
"101111000001110001110100001010100010",--15745
"111110001110001001000011100000000000",--15746
"101111000001110010000100000110011000",--15747
"111110010000000001100011000000000000",--15748
"111110001100011000000011000000000000",--15749
"111110001110001001100011000000000000",--15750
"101111000001110001110100001010000000",--15751
"111110001110001001000011100000000000",--15752
"101111000001110010000100000110001000",--15753
"111110010000000001100011000000000000",--15754
"111110001100011000000011000000000000",--15755
"111110001110001001100011000000000000",--15756
"101111000001110001110100001001000100",--15757
"111110001110001001000011100000000000",--15758
"101111000001110010000100000101110000",--15759
"111110010000000001100011000000000000",--15760
"111110001100011000000011000000000000",--15761
"111110001110001001100011000000000000",--15762
"101111000001110001110100001000010000",--15763
"111110001110001001000011100000000000",--15764
"101111000001110010000100000101010000",--15765
"111110010000000001100011000000000000",--15766
"111110001100011000000011000000000000",--15767
"111110001110001001100011000000000000",--15768
"101111000001110001110100000111001000",--15769
"111110001110001001000011100000000000",--15770
"101111000001110010000100000100110000",--15771
"111110010000000001100011000000000000",--15772
"111110001100011000000011000000000000",--15773
"111110001110001001100011000000000000",--15774
"101111000001110001110100000110000000",--15775
"111110001110001001000011100000000000",--15776
"101111000001110010000100000100010000",--15777
"111110010000000001100011000000000000",--15778
"111110001100011000000011000000000000",--15779
"111110001110001001100011000000000000",--15780
"101111000001110001110100000100010000",--15781
"111110001110001001000011100000000000",--15782
"101111000001110010000100000011100000",--15783
"111110010000000001100011000000000000",--15784
"111110001100011000000011000000000000",--15785
"111110001110001001100011000000000000",--15786
"101111000001110001110100000010000000",--15787
"111110001110001001000011100000000000",--15788
"101111000001110010000100000010100000",--15789
"111110010000000001100011000000000000",--15790
"111110001100011000000011000000000000",--15791
"111110001110001001100011000000000000",--15792
"101111000001110001110100000001000000",--15793
"111110001110000001100011000000000000",--15794
"111110001100011000000011000000000000",--15795
"111110001000001001100010000000000000",--15796
"111110001000000000010010000000000000",--15797
"111110001000011000000010000000000000",--15798
"111110000110001001000001100000000000",--15799
"010100001001000000000000000000000100",--15800
"101111001001110001000011111111001001",--15801
"101111001001100001000000111111011010",--15802
"111110001000010000110001100000000000",--15803
"000101000000000000000011110111000001",--15804
"011000001001000000000000000000000011",--15805
"101111001001110001001011111111001001",--15806
"101111001001100001000000111111011010",--15807
"111110001000010000110001100000000000",--15808
"101111000001110001000100000111110000",--15809
"111110000110001001000001100000000000",--15810
"101111001001110001000011111010100010",--15811
"101111001001100001001111100110000010",--15812
"111110000110001001000001100000000000",--15813
"101110000110110000000010000000000000",--15814
"111110000110010001000001100000000000",--15815
"101110001011111000000010000000000001",--15816
"101111001101110001100011100011010001",--15817
"101111001101100001101011011100010111",--15818
"010110001101000001000000000000000010",--15819
"101111000001110001000100000101110000",--15820
"000101000000000000000011111000110000",--15821
"001111000000000001000000000100101011",--15822
"001111000100000001100000000000000001",--15823
"111110001000010001100010000000000000",--15824
"001111000110000001100000000000000001",--15825
"111110001100100000000011000000000000",--15826
"111110001000001001100010000000000000",--15827
"111110001010011000000010100000000000",--15828
"111110001000001001010010000000000001",--15829
"010110001001000000010000000000000010",--15830
"101001000000000000100000000000000001",--15831
"000101000000000000000011110111011110",--15832
"011010001001000000100000000000000010",--15833
"101001000000000000101111111111111111",--15834
"000101000000000000000011110111011110",--15835
"101000000001111000000001000000000000",--15836
"000101000000000000000011110111011111",--15837
"111110001000011000000010000000000000",--15838
"111110001000001001000010100000000000",--15839
"101111000001110001100100001011110010",--15840
"111110001100001001010011000000000000",--15841
"101111001111110001110011110100110010",--15842
"101111001111100001110001011001000011",--15843
"111110001100001001110011000000000000",--15844
"101111000001110001110100001011001000",--15845
"111110001110001001010011100000000000",--15846
"101111000001110010000100000110101000",--15847
"111110010000000001100011000000000000",--15848
"111110001100011000000011000000000000",--15849
"111110001110001001100011000000000000",--15850
"101111000001110001110100001010100010",--15851
"111110001110001001010011100000000000",--15852
"101111000001110010000100000110011000",--15853
"111110010000000001100011000000000000",--15854
"111110001100011000000011000000000000",--15855
"111110001110001001100011000000000000",--15856
"101111000001110001110100001010000000",--15857
"111110001110001001010011100000000000",--15858
"101111000001110010000100000110001000",--15859
"111110010000000001100011000000000000",--15860
"111110001100011000000011000000000000",--15861
"111110001110001001100011000000000000",--15862
"101111000001110001110100001001000100",--15863
"111110001110001001010011100000000000",--15864
"101111000001110010000100000101110000",--15865
"111110010000000001100011000000000000",--15866
"111110001100011000000011000000000000",--15867
"111110001110001001100011000000000000",--15868
"101111000001110001110100001000010000",--15869
"111110001110001001010011100000000000",--15870
"101111000001110010000100000101010000",--15871
"111110010000000001100011000000000000",--15872
"111110001100011000000011000000000000",--15873
"111110001110001001100011000000000000",--15874
"101111000001110001110100000111001000",--15875
"111110001110001001010011100000000000",--15876
"101111000001110010000100000100110000",--15877
"111110010000000001100011000000000000",--15878
"111110001100011000000011000000000000",--15879
"111110001110001001100011000000000000",--15880
"101111000001110001110100000110000000",--15881
"111110001110001001010011100000000000",--15882
"101111000001110010000100000100010000",--15883
"111110010000000001100011000000000000",--15884
"111110001100011000000011000000000000",--15885
"111110001110001001100011000000000000",--15886
"101111000001110001110100000100010000",--15887
"111110001110001001010011100000000000",--15888
"101111000001110010000100000011100000",--15889
"111110010000000001100011000000000000",--15890
"111110001100011000000011000000000000",--15891
"111110001110001001100011000000000000",--15892
"101111000001110001110100000010000000",--15893
"111110001110001001010011100000000000",--15894
"101111000001110010000100000010100000",--15895
"111110010000000001100011000000000000",--15896
"111110001100011000000011000000000000",--15897
"111110001110001001100011000000000000",--15898
"101111000001110001110100000001000000",--15899
"111110001110000001100011000000000000",--15900
"111110001100011000000011000000000000",--15901
"111110001010001001100010100000000000",--15902
"111110001010000000010010100000000000",--15903
"111110001010011000000010100000000000",--15904
"111110001000001001010010000000000000",--15905
"010100000101000000000000000000000100",--15906
"101111001011110001010011111111001001",--15907
"101111001011100001010000111111011010",--15908
"111110001010010001000010000000000000",--15909
"000101000000000000000011111000101011",--15910
"011000000101000000000000000000000011",--15911
"101111001011110001011011111111001001",--15912
"101111001011100001010000111111011010",--15913
"111110001010010001000010000000000000",--15914
"101111000001110001010100000111110000",--15915
"111110001000001001010010000000000000",--15916
"101111001011110001010011111010100010",--15917
"101111001011100001011111100110000010",--15918
"111110001000001001010010000000000000",--15919
"101110001000110000000010100000000000",--15920
"111110001000010001010010000000000000",--15921
"101111001011110001010011111000011001",--15922
"101111001011100001011001100110011010",--15923
"101111000001110001100011111100000000",--15924
"111110001100010000110001100000000000",--15925
"111110000110001000110001100000000000",--15926
"111110001010010000110001100000000000",--15927
"101111000001110001010011111100000000",--15928
"111110001010010001000010000000000000",--15929
"111110001000001001000010000000000000",--15930
"111110000110010001000001100000000000",--15931
"011010000111000000000000000000000001",--15932
"101110000001111000000001100000000000",--15933
"101111000001110001000100001101111111",--15934
"111110001000001000110001100000000000",--15935
"101111001001110001000100000001010101",--15936
"101111001001100001000101010101010101",--15937
"111110000110001001000001100000000000",--15938
"001011000000000000110000000100100101",--15939
"001101000000000000100000000100110000",--15940
"001101000100000000010000000000000000",--15941
"001101000010000000110000000000000000",--15942
"010011000111000000000000001001101110",--15943
"001001111100000000011111111111111101",--15944
"001001111100000000101111111111111100",--15945
"010011000111011000110000000101111111",--15946
"001101000110000001000000000101101101",--15947
"001111000000000000110000000100101010",--15948
"001101001000000001010000000000000101",--15949
"001111001010000001000000000000000000",--15950
"111110000110010001000001100000000000",--15951
"001111000000000001000000000100101011",--15952
"001111001010000001010000000000000001",--15953
"111110001000010001010010000000000000",--15954
"001111000000000001010000000100101100",--15955
"001111001010000001100000000000000010",--15956
"111110001010010001100010100000000000",--15957
"001101000110000000110000000010111110",--15958
"001101001000000001010000000000000001",--15959
"011111001011000000010000000000110111",--15960
"001111000110000001100000000000000000",--15961
"111110001100010000110011000000000000",--15962
"001111000110000001110000000000000001",--15963
"111110001100001001110011000000000000",--15964
"001111000000000001110000000011111011",--15965
"111110001100001001110011100000000000",--15966
"111110001110000001000011100000000001",--15967
"001101001000000001000000000000000100",--15968
"001111001000000010000000000000000001",--15969
"010110010001000001110000000000000111",--15970
"001111000000000001110000000011111100",--15971
"111110001100001001110011100000000000",--15972
"111110001110000001010011100000000001",--15973
"001111001000000010000000000000000010",--15974
"010110010001000001110000000000000010",--15975
"001111000110000001110000000000000001",--15976
"011110001111000000000000000000100100",--15977
"001111000110000001100000000000000010",--15978
"111110001100010001000011000000000000",--15979
"001111000110000001110000000000000011",--15980
"111110001100001001110011000000000000",--15981
"001111000000000001110000000011111010",--15982
"111110001100001001110011100000000000",--15983
"111110001110000000110011100000000001",--15984
"001111001000000010000000000000000000",--15985
"010110010001000001110000000000000111",--15986
"001111000000000001110000000011111100",--15987
"111110001100001001110011100000000000",--15988
"111110001110000001010011100000000001",--15989
"001111001000000010000000000000000010",--15990
"010110010001000001110000000000000010",--15991
"001111000110000001110000000000000011",--15992
"011110001111000000000000000000010010",--15993
"001111000110000001100000000000000100",--15994
"111110001100010001010010100000000000",--15995
"001111000110000001100000000000000101",--15996
"111110001010001001100010100000000000",--15997
"001111000000000001100000000011111010",--15998
"111110001010001001100011000000000000",--15999
"111110001100000000110001100000000001",--16000
"001111001000000001100000000000000000",--16001
"010110001101000000110000000100111110",--16002
"001111000000000000110000000011111011",--16003
"111110001010001000110001100000000000",--16004
"111110000110000001000001100000000001",--16005
"001111001000000001000000000000000001",--16006
"010110001001000000110000000100111001",--16007
"001111000110000000110000000000000101",--16008
"010010000111000000000000000100110111",--16009
"001011000000000001010000000100101111",--16010
"000101000000000000000011111011011000",--16011
"001011000000000001100000000100101111",--16012
"000101000000000000000011111011011000",--16013
"001011000000000001100000000100101111",--16014
"000101000000000000000011111011011000",--16015
"011111001011000000100000000000001100",--16016
"001111000110000001100000000000000000",--16017
"011010001101000000000000000100101110",--16018
"001111000110000001100000000000000001",--16019
"111110001100001000110001100000000000",--16020
"001111000110000001100000000000000010",--16021
"111110001100001001000010000000000000",--16022
"111110000110000001000001100000000000",--16023
"001111000110000001000000000000000011",--16024
"111110001000001001010010000000000000",--16025
"111110000110000001000001100000000000",--16026
"001011000000000000110000000100101111",--16027
"000101000000000000000011111011011000",--16028
"001111000110000001100000000000000000",--16029
"010010001101000000000000000100100010",--16030
"001111000110000001110000000000000001",--16031
"111110001110001000110011100000000000",--16032
"001111000110000010000000000000000010",--16033
"111110010000001001000100000000000000",--16034
"111110001110000010000011100000000000",--16035
"001111000110000010000000000000000011",--16036
"111110010000001001010100000000000000",--16037
"111110001110000010000011100000000000",--16038
"111110000110001000110100000000000000",--16039
"001101001000000001100000000000000100",--16040
"001111001100000010010000000000000000",--16041
"111110010000001010010100000000000000",--16042
"111110001000001001000100100000000000",--16043
"001111001100000010100000000000000001",--16044
"111110010010001010100100100000000000",--16045
"111110010000000010010100000000000000",--16046
"111110001010001001010100100000000000",--16047
"001111001100000010100000000000000010",--16048
"111110010010001010100100100000000000",--16049
"111110010000000010010100000000000000",--16050
"001101001000000001100000000000000011",--16051
"011100001101000000000000000000000011",--16052
"101110010001111000000001100000000000",--16053
"011111001011000000110000000000010000",--16054
"000101000000000000000011111011000110",--16055
"111110001000001001010100100000000000",--16056
"001101001000000001100000000000001001",--16057
"001111001100000010100000000000000000",--16058
"111110010010001010100100100000000000",--16059
"111110010000000010010100000000000000",--16060
"111110001010001000110010100000000000",--16061
"001111001100000010010000000000000001",--16062
"111110001010001010010010100000000000",--16063
"111110010000000001010010100000000000",--16064
"111110000110001001000001100000000000",--16065
"001111001100000001000000000000000010",--16066
"111110000110001001000001100000000000",--16067
"111110001010000000110001100000000000",--16068
"011111001011000000110000000000000001",--16069
"111110000110010000010001100000000000",--16070
"111110001110001001110010000000000000",--16071
"111110001100001000110001100000000000",--16072
"111110001000010000110001100000000000",--16073
"010110000111000000000000000011110110",--16074
"001101001000000001000000000000000110",--16075
"011100001001000000000000000000000110",--16076
"111110000110100000000001100000000000",--16077
"111110001110010000110001100000000000",--16078
"001111000110000001000000000000000100",--16079
"111110000110001001000001100000000000",--16080
"001011000000000000110000000100101111",--16081
"000101000000000000000011111011011000",--16082
"111110000110100000000001100000000000",--16083
"111110001110000000110001100000000000",--16084
"001111000110000001000000000000000100",--16085
"111110000110001001000001100000000000",--16086
"001011000000000000110000000100101111",--16087
"001111000000000000110000000100101111",--16088
"101111001001110001001011110111001100",--16089
"101111001001100001001100110011001101",--16090
"010110001001000000110000000011100101",--16091
"001101000010000000110000000000000001",--16092
"010011000111000000000000000011100011",--16093
"001101000110000000110000000100110001",--16094
"001101000110000001000000000000000000",--16095
"010011001001000000000000000011001110",--16096
"001101001000000001010000000101101101",--16097
"001111000000000000110000000100101010",--16098
"001101001010000001100000000000000101",--16099
"001111001100000001000000000000000000",--16100
"111110000110010001000001100000000000",--16101
"001111000000000001000000000100101011",--16102
"001111001100000001010000000000000001",--16103
"111110001000010001010010000000000000",--16104
"001111000000000001010000000100101100",--16105
"001111001100000001100000000000000010",--16106
"111110001010010001100010100000000000",--16107
"001101001000000001100000000010111110",--16108
"001101001010000001110000000000000001",--16109
"011111001111000000010000000000111100",--16110
"001111001100000001100000000000000000",--16111
"111110001100010000110011000000000000",--16112
"001111001100000001110000000000000001",--16113
"111110001100001001110011000000000000",--16114
"001111000000000001110000000011111011",--16115
"111110001100001001110011100000000000",--16116
"111110001110000001000011100000000001",--16117
"001101001010000001010000000000000100",--16118
"001111001010000010000000000000000001",--16119
"010110010001000001110000000000000111",--16120
"001111000000000001110000000011111100",--16121
"111110001100001001110011100000000000",--16122
"111110001110000001010011100000000001",--16123
"001111001010000010000000000000000010",--16124
"010110010001000001110000000000000010",--16125
"001111001100000001110000000000000001",--16126
"011110001111000000000000000000101000",--16127
"001111001100000001100000000000000010",--16128
"111110001100010001000011000000000000",--16129
"001111001100000001110000000000000011",--16130
"111110001100001001110011000000000000",--16131
"001111000000000001110000000011111010",--16132
"111110001100001001110011100000000000",--16133
"111110001110000000110011100000000001",--16134
"001111001010000010000000000000000000",--16135
"010110010001000001110000000000000111",--16136
"001111000000000001110000000011111100",--16137
"111110001100001001110011100000000000",--16138
"111110001110000001010011100000000001",--16139
"001111001010000010000000000000000010",--16140
"010110010001000001110000000000000010",--16141
"001111001100000001110000000000000011",--16142
"011110001111000000000000000000010101",--16143
"001111001100000001100000000000000100",--16144
"111110001100010001010010100000000000",--16145
"001111001100000001100000000000000101",--16146
"111110001010001001100010100000000000",--16147
"001111000000000001100000000011111010",--16148
"111110001010001001100011000000000000",--16149
"111110001100000000110001100000000001",--16150
"001111001010000001100000000000000000",--16151
"010110001101000000110000000000000111",--16152
"001111000000000000110000000011111011",--16153
"111110001010001000110001100000000000",--16154
"111110000110000001000001100000000001",--16155
"001111001010000001000000000000000001",--16156
"010110001001000000110000000000000010",--16157
"001111001100000000110000000000000101",--16158
"011110000111000000000000000000000010",--16159
"101000000001111000000010100000000000",--16160
"000101000000000000000011111101111011",--16161
"001011000000000001010000000100101111",--16162
"101001000000000001010000000000000011",--16163
"000101000000000000000011111101111011",--16164
"001011000000000001100000000100101111",--16165
"101001000000000001010000000000000010",--16166
"000101000000000000000011111101111011",--16167
"001011000000000001100000000100101111",--16168
"101001000000000001010000000000000001",--16169
"000101000000000000000011111101111011",--16170
"011111001111000000100000000000001111",--16171
"001111001100000001100000000000000000",--16172
"011010001101000000000000000000001011",--16173
"001111001100000001100000000000000001",--16174
"111110001100001000110001100000000000",--16175
"001111001100000001100000000000000010",--16176
"111110001100001001000010000000000000",--16177
"111110000110000001000001100000000000",--16178
"001111001100000001000000000000000011",--16179
"111110001000001001010010000000000000",--16180
"111110000110000001000001100000000000",--16181
"001011000000000000110000000100101111",--16182
"101001000000000001010000000000000001",--16183
"000101000000000000000011111101111011",--16184
"101000000001111000000010100000000000",--16185
"000101000000000000000011111101111011",--16186
"001111001100000001100000000000000000",--16187
"011110001101000000000000000000000010",--16188
"101000000001111000000010100000000000",--16189
"000101000000000000000011111101111011",--16190
"001111001100000001110000000000000001",--16191
"111110001110001000110011100000000000",--16192
"001111001100000010000000000000000010",--16193
"111110010000001001000100000000000000",--16194
"111110001110000010000011100000000000",--16195
"001111001100000010000000000000000011",--16196
"111110010000001001010100000000000000",--16197
"111110001110000010000011100000000000",--16198
"111110000110001000110100000000000000",--16199
"001101001010000010000000000000000100",--16200
"001111010000000010010000000000000000",--16201
"111110010000001010010100000000000000",--16202
"111110001000001001000100100000000000",--16203
"001111010000000010100000000000000001",--16204
"111110010010001010100100100000000000",--16205
"111110010000000010010100000000000000",--16206
"111110001010001001010100100000000000",--16207
"001111010000000010100000000000000010",--16208
"111110010010001010100100100000000000",--16209
"111110010000000010010100000000000000",--16210
"001101001010000010000000000000000011",--16211
"011100010001000000000000000000000011",--16212
"101110010001111000000001100000000000",--16213
"011111001111000000110000000000010000",--16214
"000101000000000000000011111101100110",--16215
"111110001000001001010100100000000000",--16216
"001101001010000010000000000000001001",--16217
"001111010000000010100000000000000000",--16218
"111110010010001010100100100000000000",--16219
"111110010000000010010100000000000000",--16220
"111110001010001000110010100000000000",--16221
"001111010000000010010000000000000001",--16222
"111110001010001010010010100000000000",--16223
"111110010000000001010010100000000000",--16224
"111110000110001001000001100000000000",--16225
"001111010000000001000000000000000010",--16226
"111110000110001001000001100000000000",--16227
"111110001010000000110001100000000000",--16228
"011111001111000000110000000000000001",--16229
"111110000110010000010001100000000000",--16230
"111110001110001001110010000000000000",--16231
"111110001100001000110001100000000000",--16232
"111110001000010000110001100000000000",--16233
"010110000111000000000000000000001111",--16234
"001101001010000001010000000000000110",--16235
"011100001011000000000000000000000110",--16236
"111110000110100000000001100000000000",--16237
"111110001110010000110001100000000000",--16238
"001111001100000001000000000000000100",--16239
"111110000110001001000001100000000000",--16240
"001011000000000000110000000100101111",--16241
"000101000000000000000011111101111000",--16242
"111110000110100000000001100000000000",--16243
"111110001110000000110001100000000000",--16244
"001111001100000001000000000000000100",--16245
"111110000110001001000001100000000000",--16246
"001011000000000000110000000100101111",--16247
"101001000000000001010000000000000001",--16248
"000101000000000000000011111101111011",--16249
"101000000001111000000010100000000000",--16250
"001111000000000000110000000100101111",--16251
"010000001011000000000000000000100111",--16252
"101111001001110001001011111001001100",--16253
"101111001001100001001100110011001101",--16254
"010110001001000000110000000000100100",--16255
"101111001001110001000011110000100011",--16256
"101111001001100001001101011100001010",--16257
"111110000110000001000001100000000000",--16258
"001111000000000001000000000101100100",--16259
"111110001000001000110010000000000000",--16260
"001111000000000001010000000100101010",--16261
"111110001000000001010010000000000000",--16262
"001111000000000001010000000101100101",--16263
"111110001010001000110010100000000000",--16264
"001111000000000001100000000100101011",--16265
"111110001010000001100010100000000000",--16266
"001111000000000001100000000101100110",--16267
"111110001100001000110001100000000000",--16268
"001111000000000001100000000100101100",--16269
"111110000110000001100001100000000000",--16270
"001001111100000000111111111111111011",--16271
"101000000111111000000001000000000000",--16272
"101000000001111000000000100000000000",--16273
"101110001011111000001111100000000000",--16274
"101110000111111000000010100000000000",--16275
"101110001001111000000001100000000000",--16276
"101110111111111000000010000000000000",--16277
"001001111100000111111111111111111010",--16278
"101001111100010111100000000000000111",--16279
"000111000000000000000000011110001000",--16280
"101001111100000111100000000000000111",--16281
"001101111100000111111111111111111010",--16282
"011100000011000000000000000000101110",--16283
"101001000000000000010000000000000001",--16284
"001101111100000000101111111111111011",--16285
"101001111100010111100000000000000111",--16286
"000111000000000000000000100011100001",--16287
"101001111100000111100000000000000111",--16288
"001101111100000111111111111111111010",--16289
"011100000011000000000000000000100111",--16290
"000101000000000000000011111110101111",--16291
"001101001000000001000000000101101101",--16292
"001101001000000001000000000000000110",--16293
"010000001001000000000000000000001000",--16294
"101000000111111000000001000000000000",--16295
"101001000000000000010000000000000001",--16296
"001001111100000111111111111111111011",--16297
"101001111100010111100000000000000110",--16298
"000111000000000000000000100011100001",--16299
"101001111100000111100000000000000110",--16300
"001101111100000111111111111111111011",--16301
"011100000011000000000000000000011011",--16302
"001101111100000000011111111111111101",--16303
"001101000010000000100000000000000010",--16304
"010011000101000000000000000000001111",--16305
"001101000100000000100000000100110001",--16306
"101000000001111000000000100000000000",--16307
"001001111100000111111111111111111011",--16308
"101001111100010111100000000000000110",--16309
"000111000000000000000000100011100001",--16310
"101001111100000111100000000000000110",--16311
"001101111100000111111111111111111011",--16312
"011100000011000000000000000000010000",--16313
"101001000000000000010000000000000011",--16314
"001101111100000000101111111111111101",--16315
"101001111100010111100000000000000110",--16316
"000111000000000000000000110101111110",--16317
"101001111100000111100000000000000110",--16318
"001101111100000111111111111111111011",--16319
"011100000011000000000000000000001001",--16320
"101001000000000000010000000000000001",--16321
"001101111100000000101111111111111100",--16322
"001001111100000111111111111111111011",--16323
"101001111100010111100000000000000110",--16324
"000111000000000000000000111111111011",--16325
"101001111100000111100000000000000110",--16326
"001101111100000111111111111111111011",--16327
"011100000010000000001111100000000000",--16328
"000101000000000000000100000010110110",--16329
"001101111100000000011111111111111101",--16330
"001101000010000000100000000000000001",--16331
"010011000101000000000000000011100001",--16332
"001101000100000000100000000100110001",--16333
"001101000100000000110000000000000000",--16334
"010011000111000000000000000011001100",--16335
"001101000110000001000000000101101101",--16336
"001111000000000000110000000100101010",--16337
"001101001000000001010000000000000101",--16338
"001111001010000001000000000000000000",--16339
"111110000110010001000001100000000000",--16340
"001111000000000001000000000100101011",--16341
"001111001010000001010000000000000001",--16342
"111110001000010001010010000000000000",--16343
"001111000000000001010000000100101100",--16344
"001111001010000001100000000000000010",--16345
"111110001010010001100010100000000000",--16346
"001101000110000001010000000010111110",--16347
"001101001000000001100000000000000001",--16348
"011111001101000000010000000000111100",--16349
"001111001010000001100000000000000000",--16350
"111110001100010000110011000000000000",--16351
"001111001010000001110000000000000001",--16352
"111110001100001001110011000000000000",--16353
"001111000000000001110000000011111011",--16354
"111110001100001001110011100000000000",--16355
"111110001110000001000011100000000001",--16356
"001101001000000001000000000000000100",--16357
"001111001000000010000000000000000001",--16358
"010110010001000001110000000000000111",--16359
"001111000000000001110000000011111100",--16360
"111110001100001001110011100000000000",--16361
"111110001110000001010011100000000001",--16362
"001111001000000010000000000000000010",--16363
"010110010001000001110000000000000010",--16364
"001111001010000001110000000000000001",--16365
"011110001111000000000000000000101000",--16366
"001111001010000001100000000000000010",--16367
"111110001100010001000011000000000000",--16368
"001111001010000001110000000000000011",--16369
"111110001100001001110011000000000000",--16370
"001111000000000001110000000011111010",--16371
"111110001100001001110011100000000000",--16372
"111110001110000000110011100000000001",--16373
"001111001000000010000000000000000000",--16374
"010110010001000001110000000000000111",--16375
"001111000000000001110000000011111100",--16376
"111110001100001001110011100000000000",--16377
"111110001110000001010011100000000001",--16378
"001111001000000010000000000000000010",--16379
"010110010001000001110000000000000010",--16380
"001111001010000001110000000000000011",--16381
"011110001111000000000000000000010101",--16382
"001111001010000001100000000000000100",--16383
"111110001100010001010010100000000000",--16384
"001111001010000001100000000000000101",--16385
"111110001010001001100010100000000000",--16386
"001111000000000001100000000011111010",--16387
"111110001010001001100011000000000000",--16388
"111110001100000000110001100000000001",--16389
"001111001000000001100000000000000000",--16390
"010110001101000000110000000000000111",--16391
"001111000000000000110000000011111011",--16392
"111110001010001000110001100000000000",--16393
"111110000110000001000001100000000001",--16394
"001111001000000001000000000000000001",--16395
"010110001001000000110000000000000010",--16396
"001111001010000000110000000000000101",--16397
"011110000111000000000000000000000010",--16398
"101000000001111000000010000000000000",--16399
"000101000000000000000100000001101010",--16400
"001011000000000001010000000100101111",--16401
"101001000000000001000000000000000011",--16402
"000101000000000000000100000001101010",--16403
"001011000000000001100000000100101111",--16404
"101001000000000001000000000000000010",--16405
"000101000000000000000100000001101010",--16406
"001011000000000001100000000100101111",--16407
"101001000000000001000000000000000001",--16408
"000101000000000000000100000001101010",--16409
"011111001101000000100000000000001111",--16410
"001111001010000001100000000000000000",--16411
"011010001101000000000000000000001011",--16412
"001111001010000001100000000000000001",--16413
"111110001100001000110001100000000000",--16414
"001111001010000001100000000000000010",--16415
"111110001100001001000010000000000000",--16416
"111110000110000001000001100000000000",--16417
"001111001010000001000000000000000011",--16418
"111110001000001001010010000000000000",--16419
"111110000110000001000001100000000000",--16420
"001011000000000000110000000100101111",--16421
"101001000000000001000000000000000001",--16422
"000101000000000000000100000001101010",--16423
"101000000001111000000010000000000000",--16424
"000101000000000000000100000001101010",--16425
"001111001010000001100000000000000000",--16426
"011110001101000000000000000000000010",--16427
"101000000001111000000010000000000000",--16428
"000101000000000000000100000001101010",--16429
"001111001010000001110000000000000001",--16430
"111110001110001000110011100000000000",--16431
"001111001010000010000000000000000010",--16432
"111110010000001001000100000000000000",--16433
"111110001110000010000011100000000000",--16434
"001111001010000010000000000000000011",--16435
"111110010000001001010100000000000000",--16436
"111110001110000010000011100000000000",--16437
"111110000110001000110100000000000000",--16438
"001101001000000001110000000000000100",--16439
"001111001110000010010000000000000000",--16440
"111110010000001010010100000000000000",--16441
"111110001000001001000100100000000000",--16442
"001111001110000010100000000000000001",--16443
"111110010010001010100100100000000000",--16444
"111110010000000010010100000000000000",--16445
"111110001010001001010100100000000000",--16446
"001111001110000010100000000000000010",--16447
"111110010010001010100100100000000000",--16448
"111110010000000010010100000000000000",--16449
"001101001000000001110000000000000011",--16450
"011100001111000000000000000000000011",--16451
"101110010001111000000001100000000000",--16452
"011111001101000000110000000000010000",--16453
"000101000000000000000100000001010101",--16454
"111110001000001001010100100000000000",--16455
"001101001000000001110000000000001001",--16456
"001111001110000010100000000000000000",--16457
"111110010010001010100100100000000000",--16458
"111110010000000010010100000000000000",--16459
"111110001010001000110010100000000000",--16460
"001111001110000010010000000000000001",--16461
"111110001010001010010010100000000000",--16462
"111110010000000001010010100000000000",--16463
"111110000110001001000001100000000000",--16464
"001111001110000001000000000000000010",--16465
"111110000110001001000001100000000000",--16466
"111110001010000000110001100000000000",--16467
"011111001101000000110000000000000001",--16468
"111110000110010000010001100000000000",--16469
"111110001110001001110010000000000000",--16470
"111110001100001000110001100000000000",--16471
"111110001000010000110001100000000000",--16472
"010110000111000000000000000000001111",--16473
"001101001000000001000000000000000110",--16474
"011100001001000000000000000000000110",--16475
"111110000110100000000001100000000000",--16476
"111110001110010000110001100000000000",--16477
"001111001010000001000000000000000100",--16478
"111110000110001001000001100000000000",--16479
"001011000000000000110000000100101111",--16480
"000101000000000000000100000001100111",--16481
"111110000110100000000001100000000000",--16482
"111110001110000000110001100000000000",--16483
"001111001010000001000000000000000100",--16484
"111110000110001001000001100000000000",--16485
"001011000000000000110000000100101111",--16486
"101001000000000001000000000000000001",--16487
"000101000000000000000100000001101010",--16488
"101000000001111000000010000000000000",--16489
"001111000000000000110000000100101111",--16490
"010000001001000000000000000000100110",--16491
"101111001001110001001011111001001100",--16492
"101111001001100001001100110011001101",--16493
"010110001001000000110000000000100011",--16494
"101111001001110001000011110000100011",--16495
"101111001001100001001101011100001010",--16496
"111110000110000001000001100000000000",--16497
"001111000000000001000000000101100100",--16498
"111110001000001000110010000000000000",--16499
"001111000000000001010000000100101010",--16500
"111110001000000001010010000000000000",--16501
"001111000000000001010000000101100101",--16502
"111110001010001000110010100000000000",--16503
"001111000000000001100000000100101011",--16504
"111110001010000001100010100000000000",--16505
"001111000000000001100000000101100110",--16506
"111110001100001000110001100000000000",--16507
"001111000000000001100000000100101100",--16508
"111110000110000001100001100000000000",--16509
"001001111100000000101111111111111011",--16510
"101000000001111000000000100000000000",--16511
"101110001011111000001111100000000000",--16512
"101110000111111000000010100000000000",--16513
"101110001001111000000001100000000000",--16514
"101110111111111000000010000000000000",--16515
"001001111100000111111111111111111010",--16516
"101001111100010111100000000000000111",--16517
"000111000000000000000000011110001000",--16518
"101001111100000111100000000000000111",--16519
"001101111100000111111111111111111010",--16520
"011100000010000000001111100000000000",--16521
"101001000000000000010000000000000001",--16522
"001101111100000000101111111111111011",--16523
"101001111100010111100000000000000111",--16524
"000111000000000000000000100011100001",--16525
"101001111100000111100000000000000111",--16526
"001101111100000111111111111111111010",--16527
"011100000010000000001111100000000000",--16528
"000101000000000000000100000010011100",--16529
"001101000110000000110000000101101101",--16530
"001101000110000000110000000000000110",--16531
"010000000111000000000000000000000111",--16532
"101001000000000000010000000000000001",--16533
"001001111100000111111111111111111011",--16534
"101001111100010111100000000000000110",--16535
"000111000000000000000000100011100001",--16536
"101001111100000111100000000000000110",--16537
"001101111100000111111111111111111011",--16538
"011100000010000000001111100000000000",--16539
"001101111100000000011111111111111101",--16540
"001101000010000000100000000000000010",--16541
"010011000101000000000000000000001111",--16542
"001101000100000000100000000100110001",--16543
"101000000001111000000000100000000000",--16544
"001001111100000111111111111111111011",--16545
"101001111100010111100000000000000110",--16546
"000111000000000000000000100011100001",--16547
"101001111100000111100000000000000110",--16548
"001101111100000111111111111111111011",--16549
"011100000010000000001111100000000000",--16550
"101001000000000000010000000000000011",--16551
"001101111100000000101111111111111101",--16552
"101001111100010111100000000000000110",--16553
"000111000000000000000000110101111110",--16554
"101001111100000111100000000000000110",--16555
"001101111100000111111111111111111011",--16556
"011100000010000000001111100000000000",--16557
"101001000000000000010000000000000001",--16558
"001101111100000000101111111111111100",--16559
"001001111100000111111111111111111011",--16560
"101001111100010111100000000000000110",--16561
"000111000000000000000000111111111011",--16562
"101001111100000111100000000000000110",--16563
"001101111100000111111111111111111011",--16564
"011100000010000000001111100000000000",--16565
"001111000000000000110000000100100110",--16566
"001111000000000001000000000101100100",--16567
"111110000110001001000001100000000000",--16568
"001111000000000001000000000100100111",--16569
"001111000000000001010000000101100101",--16570
"111110001000001001010010000000000000",--16571
"111110000110000001000001100000000000",--16572
"001111000000000001000000000100101000",--16573
"001111000000000001010000000101100110",--16574
"111110001000001001010010000000000000",--16575
"111110000110000001000001100000000010",--16576
"010110000111000000000000000000000001",--16577
"000101000000000000000100000011000100",--16578
"101110000001111000000001100000000000",--16579
"001111111100000001000000000000000000",--16580
"111110001000001000110001100000000000",--16581
"001101111100000000011111111111111110",--16582
"001101000010000000010000000000000111",--16583
"001111000010000001000000000000000000",--16584
"111110000110001001000001100000000000",--16585
"001111000000000001000000000100100000",--16586
"001111000000000001010000000100100011",--16587
"111110000110001001010010100000000000",--16588
"111110001000000001010010000000000000",--16589
"001011000000000001000000000100100000",--16590
"001111000000000001000000000100100001",--16591
"001111000000000001010000000100100100",--16592
"111110000110001001010010100000000000",--16593
"111110001000000001010010000000000000",--16594
"001011000000000001000000000100100001",--16595
"001111000000000001000000000100100010",--16596
"001111000000000001010000000100100101",--16597
"111110000110001001010001100000000000",--16598
"111110001000000000110001100000000000",--16599
"001011000000000000110000000100100010",--16600
"000100000000000000001111100000000000",--16601
"010111001000000000001111100000000000",--16602
"001100000010000001000010100000000000",--16603
"001101001010000001010000000000000000",--16604
"001111001010000000110000000000000000",--16605
"001111000100000001000000000000000000",--16606
"111110000110001001000001100000000000",--16607
"001111001010000001000000000000000001",--16608
"001111000100000001010000000000000001",--16609
"111110001000001001010010000000000000",--16610
"111110000110000001000001100000000000",--16611
"001111001010000001000000000000000010",--16612
"001111000100000001010000000000000010",--16613
"111110001000001001010010000000000000",--16614
"111110000110000001000001100000000000",--16615
"001001111100000000110000000000000000",--16616
"001001111100000000101111111111111111",--16617
"001001111100000000011111111111111110",--16618
"001001111100000001001111111111111101",--16619
"011010000111000000000000001001111111",--16620
"101001001000000001010000000000000001",--16621
"001100000010000001010010100000000000",--16622
"101111001001110001000100111001101110",--16623
"101111001001100001000110101100101000",--16624
"001011000000000001000000000100101101",--16625
"001101000000000001100000000100110000",--16626
"001101001100000001110000000000000000",--16627
"001101001110000010000000000000000000",--16628
"001011111100000000111111111111111100",--16629
"001001111100000001011111111111111011",--16630
"010011010001000000000000000010000010",--16631
"001001111100000001101111111111111010",--16632
"011111010001011000110000000000001001",--16633
"101000001011111000000001100000000000",--16634
"101000001111111000000001000000000000",--16635
"101001000000000000010000000000000001",--16636
"001001111100000111111111111111111001",--16637
"101001111100010111100000000000001000",--16638
"000111000000000000000010101111001101",--16639
"101001111100000111100000000000001000",--16640
"001101111100000111111111111111111001",--16641
"000101000000000000000100000101110010",--16642
"001101010000000010010000000101101101",--16643
"001101010010000010100000000000001010",--16644
"001111010100000001000000000000000000",--16645
"001111010100000001010000000000000001",--16646
"001111010100000001100000000000000010",--16647
"001101001010000010110000000000000001",--16648
"001100010110000010000100000000000000",--16649
"001101010010000010110000000000000001",--16650
"011111010111000000010000000000111000",--16651
"001101001010000010100000000000000000",--16652
"001111010000000001110000000000000000",--16653
"111110001110010001000011100000000000",--16654
"001111010000000010000000000000000001",--16655
"111110001110001010000011100000000000",--16656
"001111010100000010000000000000000001",--16657
"111110001110001010000100000000000000",--16658
"111110010000000001010100000000000001",--16659
"001101010010000010010000000000000100",--16660
"001111010010000010010000000000000001",--16661
"010110010011000010000000000000000111",--16662
"001111010100000010000000000000000010",--16663
"111110001110001010000100000000000000",--16664
"111110010000000001100100000000000001",--16665
"001111010010000010010000000000000010",--16666
"010110010011000010000000000000000010",--16667
"001111010000000010000000000000000001",--16668
"011110010001000000000000000000100100",--16669
"001111010000000001110000000000000010",--16670
"111110001110010001010011100000000000",--16671
"001111010000000010000000000000000011",--16672
"111110001110001010000011100000000000",--16673
"001111010100000010000000000000000000",--16674
"111110001110001010000100000000000000",--16675
"111110010000000001000100000000000001",--16676
"001111010010000010010000000000000000",--16677
"010110010011000010000000000000000111",--16678
"001111010100000010000000000000000010",--16679
"111110001110001010000100000000000000",--16680
"111110010000000001100100000000000001",--16681
"001111010010000010010000000000000010",--16682
"010110010011000010000000000000000010",--16683
"001111010000000010000000000000000011",--16684
"011110010001000000000000000000010010",--16685
"001111010000000001110000000000000100",--16686
"111110001110010001100011000000000000",--16687
"001111010000000001110000000000000101",--16688
"111110001100001001110011000000000000",--16689
"001111010100000001110000000000000000",--16690
"111110001100001001110011100000000000",--16691
"111110001110000001000010000000000001",--16692
"001111010010000001110000000000000000",--16693
"010110001111000001000000000000111011",--16694
"001111010100000001000000000000000001",--16695
"111110001100001001000010000000000000",--16696
"111110001000000001010010000000000001",--16697
"001111010010000001010000000000000001",--16698
"010110001011000001000000000000110110",--16699
"001111010000000001000000000000000101",--16700
"010010001001000000000000000000110100",--16701
"001011000000000001100000000100101111",--16702
"000101000000000000000100000101100111",--16703
"001011000000000001110000000100101111",--16704
"000101000000000000000100000101100111",--16705
"001011000000000001110000000100101111",--16706
"000101000000000000000100000101100111",--16707
"011111010111000000100000000000000110",--16708
"001111010000000001000000000000000000",--16709
"011010001001000000000000000000101011",--16710
"001111010100000001010000000000000011",--16711
"111110001000001001010010000000000000",--16712
"001011000000000001000000000100101111",--16713
"000101000000000000000100000101100111",--16714
"001111010000000001110000000000000000",--16715
"010010001111000000000000000000100101",--16716
"001111010000000010000000000000000001",--16717
"111110010000001001000010000000000000",--16718
"001111010000000010000000000000000010",--16719
"111110010000001001010010100000000000",--16720
"111110001000000001010010000000000000",--16721
"001111010000000001010000000000000011",--16722
"111110001010001001100010100000000000",--16723
"111110001000000001010010000000000000",--16724
"001111010100000001010000000000000011",--16725
"111110001000001001000011000000000000",--16726
"111110001110001001010010100000000000",--16727
"111110001100010001010010100000000000",--16728
"010110001011000000000000000000011000",--16729
"001101010010000010010000000000000110",--16730
"011100010011000000000000000000000110",--16731
"111110001010100000000010100000000000",--16732
"111110001000010001010010000000000000",--16733
"001111010000000001010000000000000100",--16734
"111110001000001001010010000000000000",--16735
"001011000000000001000000000100101111",--16736
"000101000000000000000100000101100111",--16737
"111110001010100000000010100000000000",--16738
"111110001000000001010010000000000000",--16739
"001111010000000001010000000000000100",--16740
"111110001000001001010010000000000000",--16741
"001011000000000001000000000100101111",--16742
"001111000000000001000000000100101111",--16743
"001111000000000001010000000100101101",--16744
"010110001011000001000000000000001000",--16745
"101000001011111000000001100000000000",--16746
"101000001111111000000001000000000000",--16747
"101001000000000000010000000000000001",--16748
"001001111100000111111111111111111001",--16749
"101001111100010111100000000000001000",--16750
"000111000000000000000010101111001101",--16751
"101001111100000111100000000000001000",--16752
"001101111100000111111111111111111001",--16753
"101001000000000000010000000000000001",--16754
"001101111100000000101111111111111010",--16755
"001101111100000000111111111111111011",--16756
"001001111100000111111111111111111001",--16757
"101001111100010111100000000000001000",--16758
"000111000000000000000010110111111111",--16759
"101001111100000111100000000000001000",--16760
"001101111100000111111111111111111001",--16761
"001111000000000000110000000100101101",--16762
"101111001001110001001011110111001100",--16763
"101111001001100001001100110011001101",--16764
"010110000111000001000000010001101011",--16765
"101111001001110001000100110010111110",--16766
"101111001001100001001011110000100000",--16767
"010110001001000000110000010001101000",--16768
"001101000000000000010000000100101001",--16769
"001101000010000000010000000101101101",--16770
"001101000010000000100000000000000001",--16771
"011111000101000000010000000000010011",--16772
"001101111100000000101111111111111011",--16773
"001101000100000000100000000000000000",--16774
"001101000000000000110000000100101110",--16775
"001011000000000000000000000100100110",--16776
"001011000000000000000000000100100111",--16777
"001011000000000000000000000100101000",--16778
"101001000110010001000000000000000001",--16779
"101001000110010000110000000000000001",--16780
"001110000100000000110001100000000000",--16781
"011110000111000000000000000000000010",--16782
"101110000001111000000001100000000000",--16783
"000101000000000000000100000110010101",--16784
"010110000111000000000000000000000010",--16785
"101110000011111000000001100000000000",--16786
"000101000000000000000100000110010101",--16787
"101110000101111000000001100000000000",--16788
"101110000111111000000001100000000010",--16789
"001011001000000000110000000100100110",--16790
"000101000000000000000100000111101110",--16791
"011111000101000000100000000000001000",--16792
"001101000010000000100000000000000100",--16793
"001111000100010000110000000000000000",--16794
"001011000000000000110000000100100110",--16795
"001111000100010000110000000000000001",--16796
"001011000000000000110000000100100111",--16797
"001111000100010000110000000000000010",--16798
"001011000000000000110000000100101000",--16799
"000101000000000000000100000111101110",--16800
"001111000000000000110000000100101010",--16801
"001101000010000000100000000000000101",--16802
"001111000100000001000000000000000000",--16803
"111110000110010001000001100000000000",--16804
"001111000000000001000000000100101011",--16805
"001111000100000001010000000000000001",--16806
"111110001000010001010010000000000000",--16807
"001111000000000001010000000100101100",--16808
"001111000100000001100000000000000010",--16809
"111110001010010001100010100000000000",--16810
"001101000010000000100000000000000100",--16811
"001111000100000001100000000000000000",--16812
"111110000110001001100011000000000000",--16813
"001111000100000001110000000000000001",--16814
"111110001000001001110011100000000000",--16815
"001111000100000010000000000000000010",--16816
"111110001010001010000100000000000000",--16817
"001101000010000000100000000000000011",--16818
"011100000101000000000000000000000100",--16819
"001011000000000001100000000100100110",--16820
"001011000000000001110000000100100111",--16821
"001011000000000010000000000100101000",--16822
"000101000000000000000100000111010100",--16823
"001101000010000000100000000000001001",--16824
"001111000100000010010000000000000010",--16825
"111110001000001010010100100000000000",--16826
"001111000100000010100000000000000001",--16827
"111110001010001010100101000000000000",--16828
"111110010010000010100100100000000000",--16829
"101111000001110010100011111100000000",--16830
"111110010010001010100100100000000000",--16831
"111110001100000010010011000000000000",--16832
"001011000000000001100000000100100110",--16833
"001111000100000001100000000000000010",--16834
"111110000110001001100011000000000000",--16835
"001111000100000010010000000000000000",--16836
"111110001010001010010010100000000000",--16837
"111110001100000001010010100000000000",--16838
"101111000001110001100011111100000000",--16839
"111110001010001001100010100000000000",--16840
"111110001110000001010010100000000000",--16841
"001011000000000001010000000100100111",--16842
"001111000100000001010000000000000001",--16843
"111110000110001001010001100000000000",--16844
"001111000100000001010000000000000000",--16845
"111110001000001001010010000000000000",--16846
"111110000110000001000001100000000000",--16847
"101111000001110001000011111100000000",--16848
"111110000110001001000001100000000000",--16849
"111110010000000000110001100000000000",--16850
"001011000000000000110000000100101000",--16851
"001111000000000000110000000100100110",--16852
"111110000110001000110001100000000000",--16853
"001111000000000001000000000100100111",--16854
"111110001000001001000010000000000000",--16855
"111110000110000001000001100000000000",--16856
"001111000000000001000000000100101000",--16857
"111110001000001001000010000000000000",--16858
"111110000110000001000001100000000000",--16859
"111110000110100000000001100000000000",--16860
"011110000111000000000000000000000010",--16861
"101110000011111000000001100000000000",--16862
"000101000000000000000100000111100101",--16863
"001101000010000000100000000000000110",--16864
"011100000101000000000000000000000010",--16865
"111110000110011000000001100000000000",--16866
"000101000000000000000100000111100101",--16867
"111110000110011000000001100000000010",--16868
"001111000000000001000000000100100110",--16869
"111110001000001000110010000000000000",--16870
"001011000000000001000000000100100110",--16871
"001111000000000001000000000100100111",--16872
"111110001000001000110010000000000000",--16873
"001011000000000001000000000100100111",--16874
"001111000000000001000000000100101000",--16875
"111110001000001000110001100000000000",--16876
"001011000000000000110000000100101000",--16877
"001101000010000000100000000000000000",--16878
"001101000010000000110000000000001000",--16879
"001111000110000000110000000000000000",--16880
"001011000000000000110000000100100011",--16881
"001111000110000000110000000000000001",--16882
"001011000000000000110000000100100100",--16883
"001111000110000000110000000000000010",--16884
"001011000000000000110000000100100101",--16885
"001001111100000000011111111111111010",--16886
"011111000101000000010000000000100011",--16887
"001111000000000000110000000100101010",--16888
"001101000010000000100000000000000101",--16889
"001111000100000001000000000000000000",--16890
"111110000110010001000001100000000000",--16891
"101111001001110001000011110101001100",--16892
"101111001001100001001100110011001101",--16893
"111110000110001001000010000000000000",--16894
"101110001000110000000010000000000000",--16895
"101111000001110001010100000110100000",--16896
"111110001000001001010010000000000000",--16897
"111110000110010001000001100000000000",--16898
"101111000001110001000100000100100000",--16899
"001111000000000001010000000100101100",--16900
"001111000100000001100000000000000010",--16901
"111110001010010001100010100000000000",--16902
"101111001101110001100011110101001100",--16903
"101111001101100001101100110011001101",--16904
"111110001010001001100011000000000000",--16905
"101110001100110000000011000000000000",--16906
"101111000001110001110100000110100000",--16907
"111110001100001001110011000000000000",--16908
"111110001010010001100010100000000000",--16909
"101111000001110001100100000100100000",--16910
"010110001001000000110000000000000101",--16911
"010110001101000001010000000000000010",--16912
"101111000001110000110100001101111111",--16913
"000101000000000000000100001000011001",--16914
"101110000001111000000001100000000000",--16915
"000101000000000000000100001000011001",--16916
"010110001101000001010000000000000010",--16917
"101110000001111000000001100000000000",--16918
"000101000000000000000100001000011001",--16919
"101111000001110000110100001101111111",--16920
"001011000000000000110000000100100100",--16921
"000101000000000000000100001100111101",--16922
"011111000101000000100000000000001111",--16923
"001111000000000000110000000100101011",--16924
"101111000001110001000011111010000000",--16925
"111110000110001001000001100000000000",--16926
"001001111100000111111111111111111001",--16927
"000111000000000000000111011000000010",--16928
"001101111100000111111111111111111001",--16929
"111110000110001000110001100000000000",--16930
"101111000001110001000100001101111111",--16931
"111110001000001000110010000000000000",--16932
"001011000000000001000000000100100011",--16933
"101111000001110001000100001101111111",--16934
"111110000110010000010001100000000010",--16935
"111110001000001000110001100000000000",--16936
"001011000000000000110000000100100100",--16937
"000101000000000000000100001100111101",--16938
"011111000101000000110000000000011111",--16939
"001111000000000000110000000100101010",--16940
"001101000010000000100000000000000101",--16941
"001111000100000001000000000000000000",--16942
"111110000110010001000001100000000000",--16943
"001111000000000001000000000100101100",--16944
"001111000100000001010000000000000010",--16945
"111110001000010001010010000000000000",--16946
"111110000110001000110001100000000000",--16947
"111110001000001001000010000000000000",--16948
"111110000110000001000001100000000000",--16949
"111110000110100000000001100000000000",--16950
"101111001001110001000011110111001100",--16951
"101111001001100001001100110011001100",--16952
"111110000110001001000001100000000000",--16953
"101110000110110000000010000000000000",--16954
"111110000110010001000001100000000000",--16955
"101111001001110001000100000001001001",--16956
"101111001001100001000000111111011011",--16957
"111110000110001001000001100000000000",--16958
"001001111100000111111111111111111001",--16959
"000111000000000000000111010110111000",--16960
"001101111100000111111111111111111001",--16961
"111110000110001000110001100000000000",--16962
"101111000001110001000100001101111111",--16963
"111110000110001001000010000000000000",--16964
"001011000000000001000000000100100100",--16965
"111110000110010000010001100000000010",--16966
"101111000001110001000100001101111111",--16967
"111110000110001001000001100000000000",--16968
"001011000000000000110000000100100101",--16969
"000101000000000000000100001100111101",--16970
"011111000101000001000000000011110001",--16971
"001111000000000000110000000100101010",--16972
"001101000010000000100000000000000101",--16973
"001111000100000001000000000000000000",--16974
"111110000110010001000001100000000000",--16975
"001101000010000000110000000000000100",--16976
"001111000110000001000000000000000000",--16977
"111110001000100000000010000000000000",--16978
"111110000110001001000001100000000000",--16979
"001111000000000001000000000100101100",--16980
"001111000100000001010000000000000010",--16981
"111110001000010001010010000000000000",--16982
"001111000110000001010000000000000010",--16983
"111110001010100000000010100000000000",--16984
"111110001000001001010010000000000000",--16985
"111110000110001000110010100000000000",--16986
"111110001000001001000011000000000000",--16987
"111110001010000001100010100000000000",--16988
"101110000111111000000011000000000001",--16989
"101111001111110001110011100011010001",--16990
"101111001111100001111011011100010111",--16991
"010110001111000001100000000000000010",--16992
"101111000001110000110100000101110000",--16993
"000101000000000000000100001010111111",--16994
"111110000110011000000001100000000000",--16995
"111110001000001000110001100000000001",--16996
"010110000111000000010000000000000010",--16997
"101001000000000001000000000000000001",--16998
"000101000000000000000100001001101101",--16999
"011010000111000000100000000000000010",--17000
"101001000000000001001111111111111111",--17001
"000101000000000000000100001001101101",--17002
"101000000001111000000010000000000000",--17003
"000101000000000000000100001001101110",--17004
"111110000110011000000001100000000000",--17005
"111110000110001000110010000000000000",--17006
"101111000001110001100100001011110010",--17007
"111110001100001001000011000000000000",--17008
"101111001111110001110011110100110010",--17009
"101111001111100001110001011001000011",--17010
"111110001100001001110011000000000000",--17011
"101111000001110001110100001011001000",--17012
"111110001110001001000011100000000000",--17013
"101111000001110010000100000110101000",--17014
"111110010000000001100011000000000000",--17015
"111110001100011000000011000000000000",--17016
"111110001110001001100011000000000000",--17017
"101111000001110001110100001010100010",--17018
"111110001110001001000011100000000000",--17019
"101111000001110010000100000110011000",--17020
"111110010000000001100011000000000000",--17021
"111110001100011000000011000000000000",--17022
"111110001110001001100011000000000000",--17023
"101111000001110001110100001010000000",--17024
"111110001110001001000011100000000000",--17025
"101111000001110010000100000110001000",--17026
"111110010000000001100011000000000000",--17027
"111110001100011000000011000000000000",--17028
"111110001110001001100011000000000000",--17029
"101111000001110001110100001001000100",--17030
"111110001110001001000011100000000000",--17031
"101111000001110010000100000101110000",--17032
"111110010000000001100011000000000000",--17033
"111110001100011000000011000000000000",--17034
"111110001110001001100011000000000000",--17035
"101111000001110001110100001000010000",--17036
"111110001110001001000011100000000000",--17037
"101111000001110010000100000101010000",--17038
"111110010000000001100011000000000000",--17039
"111110001100011000000011000000000000",--17040
"111110001110001001100011000000000000",--17041
"101111000001110001110100000111001000",--17042
"111110001110001001000011100000000000",--17043
"101111000001110010000100000100110000",--17044
"111110010000000001100011000000000000",--17045
"111110001100011000000011000000000000",--17046
"111110001110001001100011000000000000",--17047
"101111000001110001110100000110000000",--17048
"111110001110001001000011100000000000",--17049
"101111000001110010000100000100010000",--17050
"111110010000000001100011000000000000",--17051
"111110001100011000000011000000000000",--17052
"111110001110001001100011000000000000",--17053
"101111000001110001110100000100010000",--17054
"111110001110001001000011100000000000",--17055
"101111000001110010000100000011100000",--17056
"111110010000000001100011000000000000",--17057
"111110001100011000000011000000000000",--17058
"111110001110001001100011000000000000",--17059
"101111000001110001110100000010000000",--17060
"111110001110001001000011100000000000",--17061
"101111000001110010000100000010100000",--17062
"111110010000000001100011000000000000",--17063
"111110001100011000000011000000000000",--17064
"111110001110001001100011000000000000",--17065
"101111000001110001110100000001000000",--17066
"111110001110000001100011000000000000",--17067
"111110001100011000000011000000000000",--17068
"111110001000001001100010000000000000",--17069
"111110001000000000010010000000000000",--17070
"111110001000011000000010000000000000",--17071
"111110000110001001000001100000000000",--17072
"010100001001000000000000000000000100",--17073
"101111001001110001000011111111001001",--17074
"101111001001100001000000111111011010",--17075
"111110001000010000110001100000000000",--17076
"000101000000000000000100001010111010",--17077
"011000001001000000000000000000000011",--17078
"101111001001110001001011111111001001",--17079
"101111001001100001000000111111011010",--17080
"111110001000010000110001100000000000",--17081
"101111000001110001000100000111110000",--17082
"111110000110001001000001100000000000",--17083
"101111001001110001000011111010100010",--17084
"101111001001100001001111100110000010",--17085
"111110000110001001000001100000000000",--17086
"101110000110110000000010000000000000",--17087
"111110000110010001000001100000000000",--17088
"101110001011111000000010000000000001",--17089
"101111001101110001100011100011010001",--17090
"101111001101100001101011011100010111",--17091
"010110001101000001000000000000000010",--17092
"101111000001110001000100000101110000",--17093
"000101000000000000000100001100101001",--17094
"001111000000000001000000000100101011",--17095
"001111000100000001100000000000000001",--17096
"111110001000010001100010000000000000",--17097
"001111000110000001100000000000000001",--17098
"111110001100100000000011000000000000",--17099
"111110001000001001100010000000000000",--17100
"111110001010011000000010100000000000",--17101
"111110001000001001010010000000000001",--17102
"010110001001000000010000000000000010",--17103
"101001000000000000100000000000000001",--17104
"000101000000000000000100001011010111",--17105
"011010001001000000100000000000000010",--17106
"101001000000000000101111111111111111",--17107
"000101000000000000000100001011010111",--17108
"101000000001111000000001000000000000",--17109
"000101000000000000000100001011011000",--17110
"111110001000011000000010000000000000",--17111
"111110001000001001000010100000000000",--17112
"101111000001110001100100001011110010",--17113
"111110001100001001010011000000000000",--17114
"101111001111110001110011110100110010",--17115
"101111001111100001110001011001000011",--17116
"111110001100001001110011000000000000",--17117
"101111000001110001110100001011001000",--17118
"111110001110001001010011100000000000",--17119
"101111000001110010000100000110101000",--17120
"111110010000000001100011000000000000",--17121
"111110001100011000000011000000000000",--17122
"111110001110001001100011000000000000",--17123
"101111000001110001110100001010100010",--17124
"111110001110001001010011100000000000",--17125
"101111000001110010000100000110011000",--17126
"111110010000000001100011000000000000",--17127
"111110001100011000000011000000000000",--17128
"111110001110001001100011000000000000",--17129
"101111000001110001110100001010000000",--17130
"111110001110001001010011100000000000",--17131
"101111000001110010000100000110001000",--17132
"111110010000000001100011000000000000",--17133
"111110001100011000000011000000000000",--17134
"111110001110001001100011000000000000",--17135
"101111000001110001110100001001000100",--17136
"111110001110001001010011100000000000",--17137
"101111000001110010000100000101110000",--17138
"111110010000000001100011000000000000",--17139
"111110001100011000000011000000000000",--17140
"111110001110001001100011000000000000",--17141
"101111000001110001110100001000010000",--17142
"111110001110001001010011100000000000",--17143
"101111000001110010000100000101010000",--17144
"111110010000000001100011000000000000",--17145
"111110001100011000000011000000000000",--17146
"111110001110001001100011000000000000",--17147
"101111000001110001110100000111001000",--17148
"111110001110001001010011100000000000",--17149
"101111000001110010000100000100110000",--17150
"111110010000000001100011000000000000",--17151
"111110001100011000000011000000000000",--17152
"111110001110001001100011000000000000",--17153
"101111000001110001110100000110000000",--17154
"111110001110001001010011100000000000",--17155
"101111000001110010000100000100010000",--17156
"111110010000000001100011000000000000",--17157
"111110001100011000000011000000000000",--17158
"111110001110001001100011000000000000",--17159
"101111000001110001110100000100010000",--17160
"111110001110001001010011100000000000",--17161
"101111000001110010000100000011100000",--17162
"111110010000000001100011000000000000",--17163
"111110001100011000000011000000000000",--17164
"111110001110001001100011000000000000",--17165
"101111000001110001110100000010000000",--17166
"111110001110001001010011100000000000",--17167
"101111000001110010000100000010100000",--17168
"111110010000000001100011000000000000",--17169
"111110001100011000000011000000000000",--17170
"111110001110001001100011000000000000",--17171
"101111000001110001110100000001000000",--17172
"111110001110000001100011000000000000",--17173
"111110001100011000000011000000000000",--17174
"111110001010001001100010100000000000",--17175
"111110001010000000010010100000000000",--17176
"111110001010011000000010100000000000",--17177
"111110001000001001010010000000000000",--17178
"010100000101000000000000000000000100",--17179
"101111001011110001010011111111001001",--17180
"101111001011100001010000111111011010",--17181
"111110001010010001000010000000000000",--17182
"000101000000000000000100001100100100",--17183
"011000000101000000000000000000000011",--17184
"101111001011110001011011111111001001",--17185
"101111001011100001010000111111011010",--17186
"111110001010010001000010000000000000",--17187
"101111000001110001010100000111110000",--17188
"111110001000001001010010000000000000",--17189
"101111001011110001010011111010100010",--17190
"101111001011100001011111100110000010",--17191
"111110001000001001010010000000000000",--17192
"101110001000110000000010100000000000",--17193
"111110001000010001010010000000000000",--17194
"101111001011110001010011111000011001",--17195
"101111001011100001011001100110011010",--17196
"101111000001110001100011111100000000",--17197
"111110001100010000110001100000000000",--17198
"111110000110001000110001100000000000",--17199
"111110001010010000110001100000000000",--17200
"101111000001110001010011111100000000",--17201
"111110001010010001000010000000000000",--17202
"111110001000001001000010000000000000",--17203
"111110000110010001000001100000000000",--17204
"011010000111000000000000000000000001",--17205
"101110000001111000000001100000000000",--17206
"101111000001110001000100001101111111",--17207
"111110001000001000110001100000000000",--17208
"101111001001110001000100000001010101",--17209
"101111001001100001000101010101010101",--17210
"111110000110001001000001100000000000",--17211
"001011000000000000110000000100100101",--17212
"101000000001111000000000100000000000",--17213
"001101000000000000100000000100110000",--17214
"001001111100000111111111111111111001",--17215
"101001111100010111100000000000001000",--17216
"000111000000000000000000111111111011",--17217
"101001111100000111100000000000001000",--17218
"001101111100000111111111111111111001",--17219
"011100000011000000000000001010100100",--17220
"101111000111110000111011101111011010",--17221
"101111000111100000110111010000001101",--17222
"001111111100000001001111111111111100",--17223
"111110001000001000110001100000000000",--17224
"001111000000000001000000000100100110",--17225
"001111000000000001010000000101100100",--17226
"111110001000001001010010000000000000",--17227
"001111000000000001010000000100100111",--17228
"001111000000000001100000000101100101",--17229
"111110001010001001100010100000000000",--17230
"111110001000000001010010000000000000",--17231
"001111000000000001010000000100101000",--17232
"001111000000000001100000000101100110",--17233
"111110001010001001100010100000000000",--17234
"111110001000000001010010000000000010",--17235
"010110001001000000000000000000000001",--17236
"000101000000000000000100001101010111",--17237
"101110000001111000000010000000000000",--17238
"111110000110001001000001100000000000",--17239
"001101111100000000011111111111111010",--17240
"001101000010000000010000000000000111",--17241
"001111000010000001000000000000000000",--17242
"111110000110001001000001100000000000",--17243
"001111000000000001000000000100100000",--17244
"001111000000000001010000000100100011",--17245
"111110000110001001010010100000000000",--17246
"111110001000000001010010000000000000",--17247
"001011000000000001000000000100100000",--17248
"001111000000000001000000000100100001",--17249
"001111000000000001010000000100100100",--17250
"111110000110001001010010100000000000",--17251
"111110001000000001010010000000000000",--17252
"001011000000000001000000000100100001",--17253
"001111000000000001000000000100100010",--17254
"001111000000000001010000000100100101",--17255
"111110000110001001010001100000000000",--17256
"111110001000000000110001100000000000",--17257
"001011000000000000110000000100100010",--17258
"000101000000000000000100010111101001",--17259
"001100000010000001000010100000000000",--17260
"101111001001110001000100111001101110",--17261
"101111001001100001000110101100101000",--17262
"001011000000000001000000000100101101",--17263
"001101000000000001100000000100110000",--17264
"001101001100000001110000000000000000",--17265
"001101001110000010000000000000000000",--17266
"001011111100000000111111111111111100",--17267
"001001111100000001011111111111111011",--17268
"010011010001000000000000000010000010",--17269
"001001111100000001101111111111111010",--17270
"011111010001011000110000000000001001",--17271
"101000001011111000000001100000000000",--17272
"101000001111111000000001000000000000",--17273
"101001000000000000010000000000000001",--17274
"001001111100000111111111111111111001",--17275
"101001111100010111100000000000001000",--17276
"000111000000000000000010101111001101",--17277
"101001111100000111100000000000001000",--17278
"001101111100000111111111111111111001",--17279
"000101000000000000000100001111110000",--17280
"001101010000000010010000000101101101",--17281
"001101010010000010100000000000001010",--17282
"001111010100000001000000000000000000",--17283
"001111010100000001010000000000000001",--17284
"001111010100000001100000000000000010",--17285
"001101001010000010110000000000000001",--17286
"001100010110000010000100000000000000",--17287
"001101010010000010110000000000000001",--17288
"011111010111000000010000000000111000",--17289
"001101001010000010100000000000000000",--17290
"001111010000000001110000000000000000",--17291
"111110001110010001000011100000000000",--17292
"001111010000000010000000000000000001",--17293
"111110001110001010000011100000000000",--17294
"001111010100000010000000000000000001",--17295
"111110001110001010000100000000000000",--17296
"111110010000000001010100000000000001",--17297
"001101010010000010010000000000000100",--17298
"001111010010000010010000000000000001",--17299
"010110010011000010000000000000000111",--17300
"001111010100000010000000000000000010",--17301
"111110001110001010000100000000000000",--17302
"111110010000000001100100000000000001",--17303
"001111010010000010010000000000000010",--17304
"010110010011000010000000000000000010",--17305
"001111010000000010000000000000000001",--17306
"011110010001000000000000000000100100",--17307
"001111010000000001110000000000000010",--17308
"111110001110010001010011100000000000",--17309
"001111010000000010000000000000000011",--17310
"111110001110001010000011100000000000",--17311
"001111010100000010000000000000000000",--17312
"111110001110001010000100000000000000",--17313
"111110010000000001000100000000000001",--17314
"001111010010000010010000000000000000",--17315
"010110010011000010000000000000000111",--17316
"001111010100000010000000000000000010",--17317
"111110001110001010000100000000000000",--17318
"111110010000000001100100000000000001",--17319
"001111010010000010010000000000000010",--17320
"010110010011000010000000000000000010",--17321
"001111010000000010000000000000000011",--17322
"011110010001000000000000000000010010",--17323
"001111010000000001110000000000000100",--17324
"111110001110010001100011000000000000",--17325
"001111010000000001110000000000000101",--17326
"111110001100001001110011000000000000",--17327
"001111010100000001110000000000000000",--17328
"111110001100001001110011100000000000",--17329
"111110001110000001000010000000000001",--17330
"001111010010000001110000000000000000",--17331
"010110001111000001000000000000111011",--17332
"001111010100000001000000000000000001",--17333
"111110001100001001000010000000000000",--17334
"111110001000000001010010000000000001",--17335
"001111010010000001010000000000000001",--17336
"010110001011000001000000000000110110",--17337
"001111010000000001000000000000000101",--17338
"010010001001000000000000000000110100",--17339
"001011000000000001100000000100101111",--17340
"000101000000000000000100001111100101",--17341
"001011000000000001110000000100101111",--17342
"000101000000000000000100001111100101",--17343
"001011000000000001110000000100101111",--17344
"000101000000000000000100001111100101",--17345
"011111010111000000100000000000000110",--17346
"001111010000000001000000000000000000",--17347
"011010001001000000000000000000101011",--17348
"001111010100000001010000000000000011",--17349
"111110001000001001010010000000000000",--17350
"001011000000000001000000000100101111",--17351
"000101000000000000000100001111100101",--17352
"001111010000000001110000000000000000",--17353
"010010001111000000000000000000100101",--17354
"001111010000000010000000000000000001",--17355
"111110010000001001000010000000000000",--17356
"001111010000000010000000000000000010",--17357
"111110010000001001010010100000000000",--17358
"111110001000000001010010000000000000",--17359
"001111010000000001010000000000000011",--17360
"111110001010001001100010100000000000",--17361
"111110001000000001010010000000000000",--17362
"001111010100000001010000000000000011",--17363
"111110001000001001000011000000000000",--17364
"111110001110001001010010100000000000",--17365
"111110001100010001010010100000000000",--17366
"010110001011000000000000000000011000",--17367
"001101010010000010010000000000000110",--17368
"011100010011000000000000000000000110",--17369
"111110001010100000000010100000000000",--17370
"111110001000010001010010000000000000",--17371
"001111010000000001010000000000000100",--17372
"111110001000001001010010000000000000",--17373
"001011000000000001000000000100101111",--17374
"000101000000000000000100001111100101",--17375
"111110001010100000000010100000000000",--17376
"111110001000000001010010000000000000",--17377
"001111010000000001010000000000000100",--17378
"111110001000001001010010000000000000",--17379
"001011000000000001000000000100101111",--17380
"001111000000000001000000000100101111",--17381
"001111000000000001010000000100101101",--17382
"010110001011000001000000000000001000",--17383
"101000001011111000000001100000000000",--17384
"101000001111111000000001000000000000",--17385
"101001000000000000010000000000000001",--17386
"001001111100000111111111111111111001",--17387
"101001111100010111100000000000001000",--17388
"000111000000000000000010101111001101",--17389
"101001111100000111100000000000001000",--17390
"001101111100000111111111111111111001",--17391
"101001000000000000010000000000000001",--17392
"001101111100000000101111111111111010",--17393
"001101111100000000111111111111111011",--17394
"001001111100000111111111111111111001",--17395
"101001111100010111100000000000001000",--17396
"000111000000000000000010110111111111",--17397
"101001111100000111100000000000001000",--17398
"001101111100000111111111111111111001",--17399
"001111000000000000110000000100101101",--17400
"101111001001110001001011110111001100",--17401
"101111001001100001001100110011001101",--17402
"010110000111000001000000000111101101",--17403
"101111001001110001000100110010111110",--17404
"101111001001100001001011110000100000",--17405
"010110001001000000110000000111101010",--17406
"001101000000000000010000000100101001",--17407
"001101000010000000010000000101101101",--17408
"001101000010000000100000000000000001",--17409
"011111000101000000010000000000010011",--17410
"001101111100000000101111111111111011",--17411
"001101000100000000100000000000000000",--17412
"001101000000000000110000000100101110",--17413
"001011000000000000000000000100100110",--17414
"001011000000000000000000000100100111",--17415
"001011000000000000000000000100101000",--17416
"101001000110010001000000000000000001",--17417
"101001000110010000110000000000000001",--17418
"001110000100000000110001100000000000",--17419
"011110000111000000000000000000000010",--17420
"101110000001111000000001100000000000",--17421
"000101000000000000000100010000010011",--17422
"010110000111000000000000000000000010",--17423
"101110000011111000000001100000000000",--17424
"000101000000000000000100010000010011",--17425
"101110000101111000000001100000000000",--17426
"101110000111111000000001100000000010",--17427
"001011001000000000110000000100100110",--17428
"000101000000000000000100010001101100",--17429
"011111000101000000100000000000001000",--17430
"001101000010000000100000000000000100",--17431
"001111000100010000110000000000000000",--17432
"001011000000000000110000000100100110",--17433
"001111000100010000110000000000000001",--17434
"001011000000000000110000000100100111",--17435
"001111000100010000110000000000000010",--17436
"001011000000000000110000000100101000",--17437
"000101000000000000000100010001101100",--17438
"001111000000000000110000000100101010",--17439
"001101000010000000100000000000000101",--17440
"001111000100000001000000000000000000",--17441
"111110000110010001000001100000000000",--17442
"001111000000000001000000000100101011",--17443
"001111000100000001010000000000000001",--17444
"111110001000010001010010000000000000",--17445
"001111000000000001010000000100101100",--17446
"001111000100000001100000000000000010",--17447
"111110001010010001100010100000000000",--17448
"001101000010000000100000000000000100",--17449
"001111000100000001100000000000000000",--17450
"111110000110001001100011000000000000",--17451
"001111000100000001110000000000000001",--17452
"111110001000001001110011100000000000",--17453
"001111000100000010000000000000000010",--17454
"111110001010001010000100000000000000",--17455
"001101000010000000100000000000000011",--17456
"011100000101000000000000000000000100",--17457
"001011000000000001100000000100100110",--17458
"001011000000000001110000000100100111",--17459
"001011000000000010000000000100101000",--17460
"000101000000000000000100010001010010",--17461
"001101000010000000100000000000001001",--17462
"001111000100000010010000000000000010",--17463
"111110001000001010010100100000000000",--17464
"001111000100000010100000000000000001",--17465
"111110001010001010100101000000000000",--17466
"111110010010000010100100100000000000",--17467
"101111000001110010100011111100000000",--17468
"111110010010001010100100100000000000",--17469
"111110001100000010010011000000000000",--17470
"001011000000000001100000000100100110",--17471
"001111000100000001100000000000000010",--17472
"111110000110001001100011000000000000",--17473
"001111000100000010010000000000000000",--17474
"111110001010001010010010100000000000",--17475
"111110001100000001010010100000000000",--17476
"101111000001110001100011111100000000",--17477
"111110001010001001100010100000000000",--17478
"111110001110000001010010100000000000",--17479
"001011000000000001010000000100100111",--17480
"001111000100000001010000000000000001",--17481
"111110000110001001010001100000000000",--17482
"001111000100000001010000000000000000",--17483
"111110001000001001010010000000000000",--17484
"111110000110000001000001100000000000",--17485
"101111000001110001000011111100000000",--17486
"111110000110001001000001100000000000",--17487
"111110010000000000110001100000000000",--17488
"001011000000000000110000000100101000",--17489
"001111000000000000110000000100100110",--17490
"111110000110001000110001100000000000",--17491
"001111000000000001000000000100100111",--17492
"111110001000001001000010000000000000",--17493
"111110000110000001000001100000000000",--17494
"001111000000000001000000000100101000",--17495
"111110001000001001000010000000000000",--17496
"111110000110000001000001100000000000",--17497
"111110000110100000000001100000000000",--17498
"011110000111000000000000000000000010",--17499
"101110000011111000000001100000000000",--17500
"000101000000000000000100010001100011",--17501
"001101000010000000100000000000000110",--17502
"011100000101000000000000000000000010",--17503
"111110000110011000000001100000000000",--17504
"000101000000000000000100010001100011",--17505
"111110000110011000000001100000000010",--17506
"001111000000000001000000000100100110",--17507
"111110001000001000110010000000000000",--17508
"001011000000000001000000000100100110",--17509
"001111000000000001000000000100100111",--17510
"111110001000001000110010000000000000",--17511
"001011000000000001000000000100100111",--17512
"001111000000000001000000000100101000",--17513
"111110001000001000110001100000000000",--17514
"001011000000000000110000000100101000",--17515
"001101000010000000100000000000000000",--17516
"001101000010000000110000000000001000",--17517
"001111000110000000110000000000000000",--17518
"001011000000000000110000000100100011",--17519
"001111000110000000110000000000000001",--17520
"001011000000000000110000000100100100",--17521
"001111000110000000110000000000000010",--17522
"001011000000000000110000000100100101",--17523
"001001111100000000011111111111111010",--17524
"011111000101000000010000000000100011",--17525
"001111000000000000110000000100101010",--17526
"001101000010000000100000000000000101",--17527
"001111000100000001000000000000000000",--17528
"111110000110010001000001100000000000",--17529
"101111001001110001000011110101001100",--17530
"101111001001100001001100110011001101",--17531
"111110000110001001000010000000000000",--17532
"101110001000110000000010000000000000",--17533
"101111000001110001010100000110100000",--17534
"111110001000001001010010000000000000",--17535
"111110000110010001000001100000000000",--17536
"101111000001110001000100000100100000",--17537
"001111000000000001010000000100101100",--17538
"001111000100000001100000000000000010",--17539
"111110001010010001100010100000000000",--17540
"101111001101110001100011110101001100",--17541
"101111001101100001101100110011001101",--17542
"111110001010001001100011000000000000",--17543
"101110001100110000000011000000000000",--17544
"101111000001110001110100000110100000",--17545
"111110001100001001110011000000000000",--17546
"111110001010010001100010100000000000",--17547
"101111000001110001100100000100100000",--17548
"010110001001000000110000000000000101",--17549
"010110001101000001010000000000000010",--17550
"101111000001110000110100001101111111",--17551
"000101000000000000000100010010010111",--17552
"101110000001111000000001100000000000",--17553
"000101000000000000000100010010010111",--17554
"010110001101000001010000000000000010",--17555
"101110000001111000000001100000000000",--17556
"000101000000000000000100010010010111",--17557
"101111000001110000110100001101111111",--17558
"001011000000000000110000000100100100",--17559
"000101000000000000000100010110111011",--17560
"011111000101000000100000000000001111",--17561
"001111000000000000110000000100101011",--17562
"101111000001110001000011111010000000",--17563
"111110000110001001000001100000000000",--17564
"001001111100000111111111111111111001",--17565
"000111000000000000000111011000000010",--17566
"001101111100000111111111111111111001",--17567
"111110000110001000110001100000000000",--17568
"101111000001110001000100001101111111",--17569
"111110001000001000110010000000000000",--17570
"001011000000000001000000000100100011",--17571
"101111000001110001000100001101111111",--17572
"111110000110010000010001100000000010",--17573
"111110001000001000110001100000000000",--17574
"001011000000000000110000000100100100",--17575
"000101000000000000000100010110111011",--17576
"011111000101000000110000000000011111",--17577
"001111000000000000110000000100101010",--17578
"001101000010000000100000000000000101",--17579
"001111000100000001000000000000000000",--17580
"111110000110010001000001100000000000",--17581
"001111000000000001000000000100101100",--17582
"001111000100000001010000000000000010",--17583
"111110001000010001010010000000000000",--17584
"111110000110001000110001100000000000",--17585
"111110001000001001000010000000000000",--17586
"111110000110000001000001100000000000",--17587
"111110000110100000000001100000000000",--17588
"101111001001110001000011110111001100",--17589
"101111001001100001001100110011001100",--17590
"111110000110001001000001100000000000",--17591
"101110000110110000000010000000000000",--17592
"111110000110010001000001100000000000",--17593
"101111001001110001000100000001001001",--17594
"101111001001100001000000111111011011",--17595
"111110000110001001000001100000000000",--17596
"001001111100000111111111111111111001",--17597
"000111000000000000000111010110111000",--17598
"001101111100000111111111111111111001",--17599
"111110000110001000110001100000000000",--17600
"101111000001110001000100001101111111",--17601
"111110000110001001000010000000000000",--17602
"001011000000000001000000000100100100",--17603
"111110000110010000010001100000000010",--17604
"101111000001110001000100001101111111",--17605
"111110000110001001000001100000000000",--17606
"001011000000000000110000000100100101",--17607
"000101000000000000000100010110111011",--17608
"011111000101000001000000000011110001",--17609
"001111000000000000110000000100101010",--17610
"001101000010000000100000000000000101",--17611
"001111000100000001000000000000000000",--17612
"111110000110010001000001100000000000",--17613
"001101000010000000110000000000000100",--17614
"001111000110000001000000000000000000",--17615
"111110001000100000000010000000000000",--17616
"111110000110001001000001100000000000",--17617
"001111000000000001000000000100101100",--17618
"001111000100000001010000000000000010",--17619
"111110001000010001010010000000000000",--17620
"001111000110000001010000000000000010",--17621
"111110001010100000000010100000000000",--17622
"111110001000001001010010000000000000",--17623
"111110000110001000110010100000000000",--17624
"111110001000001001000011000000000000",--17625
"111110001010000001100010100000000000",--17626
"101110000111111000000011000000000001",--17627
"101111001111110001110011100011010001",--17628
"101111001111100001111011011100010111",--17629
"010110001111000001100000000000000010",--17630
"101111000001110000110100000101110000",--17631
"000101000000000000000100010100111101",--17632
"111110000110011000000001100000000000",--17633
"111110001000001000110001100000000001",--17634
"010110000111000000010000000000000010",--17635
"101001000000000001000000000000000001",--17636
"000101000000000000000100010011101011",--17637
"011010000111000000100000000000000010",--17638
"101001000000000001001111111111111111",--17639
"000101000000000000000100010011101011",--17640
"101000000001111000000010000000000000",--17641
"000101000000000000000100010011101100",--17642
"111110000110011000000001100000000000",--17643
"111110000110001000110010000000000000",--17644
"101111000001110001100100001011110010",--17645
"111110001100001001000011000000000000",--17646
"101111001111110001110011110100110010",--17647
"101111001111100001110001011001000011",--17648
"111110001100001001110011000000000000",--17649
"101111000001110001110100001011001000",--17650
"111110001110001001000011100000000000",--17651
"101111000001110010000100000110101000",--17652
"111110010000000001100011000000000000",--17653
"111110001100011000000011000000000000",--17654
"111110001110001001100011000000000000",--17655
"101111000001110001110100001010100010",--17656
"111110001110001001000011100000000000",--17657
"101111000001110010000100000110011000",--17658
"111110010000000001100011000000000000",--17659
"111110001100011000000011000000000000",--17660
"111110001110001001100011000000000000",--17661
"101111000001110001110100001010000000",--17662
"111110001110001001000011100000000000",--17663
"101111000001110010000100000110001000",--17664
"111110010000000001100011000000000000",--17665
"111110001100011000000011000000000000",--17666
"111110001110001001100011000000000000",--17667
"101111000001110001110100001001000100",--17668
"111110001110001001000011100000000000",--17669
"101111000001110010000100000101110000",--17670
"111110010000000001100011000000000000",--17671
"111110001100011000000011000000000000",--17672
"111110001110001001100011000000000000",--17673
"101111000001110001110100001000010000",--17674
"111110001110001001000011100000000000",--17675
"101111000001110010000100000101010000",--17676
"111110010000000001100011000000000000",--17677
"111110001100011000000011000000000000",--17678
"111110001110001001100011000000000000",--17679
"101111000001110001110100000111001000",--17680
"111110001110001001000011100000000000",--17681
"101111000001110010000100000100110000",--17682
"111110010000000001100011000000000000",--17683
"111110001100011000000011000000000000",--17684
"111110001110001001100011000000000000",--17685
"101111000001110001110100000110000000",--17686
"111110001110001001000011100000000000",--17687
"101111000001110010000100000100010000",--17688
"111110010000000001100011000000000000",--17689
"111110001100011000000011000000000000",--17690
"111110001110001001100011000000000000",--17691
"101111000001110001110100000100010000",--17692
"111110001110001001000011100000000000",--17693
"101111000001110010000100000011100000",--17694
"111110010000000001100011000000000000",--17695
"111110001100011000000011000000000000",--17696
"111110001110001001100011000000000000",--17697
"101111000001110001110100000010000000",--17698
"111110001110001001000011100000000000",--17699
"101111000001110010000100000010100000",--17700
"111110010000000001100011000000000000",--17701
"111110001100011000000011000000000000",--17702
"111110001110001001100011000000000000",--17703
"101111000001110001110100000001000000",--17704
"111110001110000001100011000000000000",--17705
"111110001100011000000011000000000000",--17706
"111110001000001001100010000000000000",--17707
"111110001000000000010010000000000000",--17708
"111110001000011000000010000000000000",--17709
"111110000110001001000001100000000000",--17710
"010100001001000000000000000000000100",--17711
"101111001001110001000011111111001001",--17712
"101111001001100001000000111111011010",--17713
"111110001000010000110001100000000000",--17714
"000101000000000000000100010100111000",--17715
"011000001001000000000000000000000011",--17716
"101111001001110001001011111111001001",--17717
"101111001001100001000000111111011010",--17718
"111110001000010000110001100000000000",--17719
"101111000001110001000100000111110000",--17720
"111110000110001001000001100000000000",--17721
"101111001001110001000011111010100010",--17722
"101111001001100001001111100110000010",--17723
"111110000110001001000001100000000000",--17724
"101110000110110000000010000000000000",--17725
"111110000110010001000001100000000000",--17726
"101110001011111000000010000000000001",--17727
"101111001101110001100011100011010001",--17728
"101111001101100001101011011100010111",--17729
"010110001101000001000000000000000010",--17730
"101111000001110001000100000101110000",--17731
"000101000000000000000100010110100111",--17732
"001111000000000001000000000100101011",--17733
"001111000100000001100000000000000001",--17734
"111110001000010001100010000000000000",--17735
"001111000110000001100000000000000001",--17736
"111110001100100000000011000000000000",--17737
"111110001000001001100010000000000000",--17738
"111110001010011000000010100000000000",--17739
"111110001000001001010010000000000001",--17740
"010110001001000000010000000000000010",--17741
"101001000000000000100000000000000001",--17742
"000101000000000000000100010101010101",--17743
"011010001001000000100000000000000010",--17744
"101001000000000000101111111111111111",--17745
"000101000000000000000100010101010101",--17746
"101000000001111000000001000000000000",--17747
"000101000000000000000100010101010110",--17748
"111110001000011000000010000000000000",--17749
"111110001000001001000010100000000000",--17750
"101111000001110001100100001011110010",--17751
"111110001100001001010011000000000000",--17752
"101111001111110001110011110100110010",--17753
"101111001111100001110001011001000011",--17754
"111110001100001001110011000000000000",--17755
"101111000001110001110100001011001000",--17756
"111110001110001001010011100000000000",--17757
"101111000001110010000100000110101000",--17758
"111110010000000001100011000000000000",--17759
"111110001100011000000011000000000000",--17760
"111110001110001001100011000000000000",--17761
"101111000001110001110100001010100010",--17762
"111110001110001001010011100000000000",--17763
"101111000001110010000100000110011000",--17764
"111110010000000001100011000000000000",--17765
"111110001100011000000011000000000000",--17766
"111110001110001001100011000000000000",--17767
"101111000001110001110100001010000000",--17768
"111110001110001001010011100000000000",--17769
"101111000001110010000100000110001000",--17770
"111110010000000001100011000000000000",--17771
"111110001100011000000011000000000000",--17772
"111110001110001001100011000000000000",--17773
"101111000001110001110100001001000100",--17774
"111110001110001001010011100000000000",--17775
"101111000001110010000100000101110000",--17776
"111110010000000001100011000000000000",--17777
"111110001100011000000011000000000000",--17778
"111110001110001001100011000000000000",--17779
"101111000001110001110100001000010000",--17780
"111110001110001001010011100000000000",--17781
"101111000001110010000100000101010000",--17782
"111110010000000001100011000000000000",--17783
"111110001100011000000011000000000000",--17784
"111110001110001001100011000000000000",--17785
"101111000001110001110100000111001000",--17786
"111110001110001001010011100000000000",--17787
"101111000001110010000100000100110000",--17788
"111110010000000001100011000000000000",--17789
"111110001100011000000011000000000000",--17790
"111110001110001001100011000000000000",--17791
"101111000001110001110100000110000000",--17792
"111110001110001001010011100000000000",--17793
"101111000001110010000100000100010000",--17794
"111110010000000001100011000000000000",--17795
"111110001100011000000011000000000000",--17796
"111110001110001001100011000000000000",--17797
"101111000001110001110100000100010000",--17798
"111110001110001001010011100000000000",--17799
"101111000001110010000100000011100000",--17800
"111110010000000001100011000000000000",--17801
"111110001100011000000011000000000000",--17802
"111110001110001001100011000000000000",--17803
"101111000001110001110100000010000000",--17804
"111110001110001001010011100000000000",--17805
"101111000001110010000100000010100000",--17806
"111110010000000001100011000000000000",--17807
"111110001100011000000011000000000000",--17808
"111110001110001001100011000000000000",--17809
"101111000001110001110100000001000000",--17810
"111110001110000001100011000000000000",--17811
"111110001100011000000011000000000000",--17812
"111110001010001001100010100000000000",--17813
"111110001010000000010010100000000000",--17814
"111110001010011000000010100000000000",--17815
"111110001000001001010010000000000000",--17816
"010100000101000000000000000000000100",--17817
"101111001011110001010011111111001001",--17818
"101111001011100001010000111111011010",--17819
"111110001010010001000010000000000000",--17820
"000101000000000000000100010110100010",--17821
"011000000101000000000000000000000011",--17822
"101111001011110001011011111111001001",--17823
"101111001011100001010000111111011010",--17824
"111110001010010001000010000000000000",--17825
"101111000001110001010100000111110000",--17826
"111110001000001001010010000000000000",--17827
"101111001011110001010011111010100010",--17828
"101111001011100001011111100110000010",--17829
"111110001000001001010010000000000000",--17830
"101110001000110000000010100000000000",--17831
"111110001000010001010010000000000000",--17832
"101111001011110001010011111000011001",--17833
"101111001011100001011001100110011010",--17834
"101111000001110001100011111100000000",--17835
"111110001100010000110001100000000000",--17836
"111110000110001000110001100000000000",--17837
"111110001010010000110001100000000000",--17838
"101111000001110001010011111100000000",--17839
"111110001010010001000010000000000000",--17840
"111110001000001001000010000000000000",--17841
"111110000110010001000001100000000000",--17842
"011010000111000000000000000000000001",--17843
"101110000001111000000001100000000000",--17844
"101111000001110001000100001101111111",--17845
"111110001000001000110001100000000000",--17846
"101111001001110001000100000001010101",--17847
"101111001001100001000101010101010101",--17848
"111110000110001001000001100000000000",--17849
"001011000000000000110000000100100101",--17850
"101000000001111000000000100000000000",--17851
"001101000000000000100000000100110000",--17852
"001001111100000111111111111111111001",--17853
"101001111100010111100000000000001000",--17854
"000111000000000000000000111111111011",--17855
"101001111100000111100000000000001000",--17856
"001101111100000111111111111111111001",--17857
"011100000011000000000000000000100110",--17858
"101111000111110000110011101111011010",--17859
"101111000111100000110111010000001101",--17860
"001111111100000001001111111111111100",--17861
"111110001000001000110001100000000000",--17862
"001111000000000001000000000100100110",--17863
"001111000000000001010000000101100100",--17864
"111110001000001001010010000000000000",--17865
"001111000000000001010000000100100111",--17866
"001111000000000001100000000101100101",--17867
"111110001010001001100010100000000000",--17868
"111110001000000001010010000000000000",--17869
"001111000000000001010000000100101000",--17870
"001111000000000001100000000101100110",--17871
"111110001010001001100010100000000000",--17872
"111110001000000001010010000000000010",--17873
"010110001001000000000000000000000001",--17874
"000101000000000000000100010111010101",--17875
"101110000001111000000010000000000000",--17876
"111110000110001001000001100000000000",--17877
"001101111100000000011111111111111010",--17878
"001101000010000000010000000000000111",--17879
"001111000010000001000000000000000000",--17880
"111110000110001001000001100000000000",--17881
"001111000000000001000000000100100000",--17882
"001111000000000001010000000100100011",--17883
"111110000110001001010010100000000000",--17884
"111110001000000001010010000000000000",--17885
"001011000000000001000000000100100000",--17886
"001111000000000001000000000100100001",--17887
"001111000000000001010000000100100100",--17888
"111110000110001001010010100000000000",--17889
"111110001000000001010010000000000000",--17890
"001011000000000001000000000100100001",--17891
"001111000000000001000000000100100010",--17892
"001111000000000001010000000100100101",--17893
"111110000110001001010001100000000000",--17894
"111110001000000000110001100000000000",--17895
"001011000000000000110000000100100010",--17896
"001101111100000000011111111111111101",--17897
"101001000010010000010000000000000010",--17898
"010111000010000000001111100000000000",--17899
"001101111100000000111111111111111110",--17900
"001100000110000000010001000000000000",--17901
"001101000100000000100000000000000000",--17902
"001111000100000000110000000000000000",--17903
"001101111100000001001111111111111111",--17904
"001111001000000001000000000000000000",--17905
"111110000110001001000001100000000000",--17906
"001111000100000001000000000000000001",--17907
"001111001000000001010000000000000001",--17908
"111110001000001001010010000000000000",--17909
"111110000110000001000001100000000000",--17910
"001111000100000001000000000000000010",--17911
"001111001000000001010000000000000010",--17912
"111110001000001001010010000000000000",--17913
"111110000110000001000001100000000000",--17914
"001001111100000000011111111111111011",--17915
"011010000111000000000000001011000111",--17916
"101001000010000000100000000000000001",--17917
"001100000110000000100001100000000000",--17918
"101111001001110001000100111001101110",--17919
"101111001001100001000110101100101000",--17920
"001011000000000001000000000100101101",--17921
"001101000000000000100000000100110000",--17922
"001011111100000000111111111111111010",--17923
"001001111100000000111111111111111001",--17924
"101000000001111000000000100000000000",--17925
"001001111100000111111111111111111000",--17926
"101001111100010111100000000000001001",--17927
"000111000000000000000010110111111111",--17928
"101001111100000111100000000000001001",--17929
"001101111100000111111111111111111000",--17930
"001111000000000000110000000100101101",--17931
"101111001001110001001011110111001100",--17932
"101111001001100001001100110011001101",--17933
"010110000111000001000000010101111010",--17934
"101111001001110001000100110010111110",--17935
"101111001001100001001011110000100000",--17936
"010110001001000000110000010101110111",--17937
"001101000000000000010000000100101001",--17938
"001101000010000000010000000101101101",--17939
"001101000010000000100000000000000001",--17940
"011111000101000000010000000000010011",--17941
"001101111100000000101111111111111001",--17942
"001101000100000000100000000000000000",--17943
"001101000000000000110000000100101110",--17944
"001011000000000000000000000100100110",--17945
"001011000000000000000000000100100111",--17946
"001011000000000000000000000100101000",--17947
"101001000110010001000000000000000001",--17948
"101001000110010000110000000000000001",--17949
"001110000100000000110001100000000000",--17950
"011110000111000000000000000000000010",--17951
"101110000001111000000001100000000000",--17952
"000101000000000000000100011000100110",--17953
"010110000111000000000000000000000010",--17954
"101110000011111000000001100000000000",--17955
"000101000000000000000100011000100110",--17956
"101110000101111000000001100000000000",--17957
"101110000111111000000001100000000010",--17958
"001011001000000000110000000100100110",--17959
"000101000000000000000100011001111111",--17960
"011111000101000000100000000000001000",--17961
"001101000010000000100000000000000100",--17962
"001111000100010000110000000000000000",--17963
"001011000000000000110000000100100110",--17964
"001111000100010000110000000000000001",--17965
"001011000000000000110000000100100111",--17966
"001111000100010000110000000000000010",--17967
"001011000000000000110000000100101000",--17968
"000101000000000000000100011001111111",--17969
"001111000000000000110000000100101010",--17970
"001101000010000000100000000000000101",--17971
"001111000100000001000000000000000000",--17972
"111110000110010001000001100000000000",--17973
"001111000000000001000000000100101011",--17974
"001111000100000001010000000000000001",--17975
"111110001000010001010010000000000000",--17976
"001111000000000001010000000100101100",--17977
"001111000100000001100000000000000010",--17978
"111110001010010001100010100000000000",--17979
"001101000010000000100000000000000100",--17980
"001111000100000001100000000000000000",--17981
"111110000110001001100011000000000000",--17982
"001111000100000001110000000000000001",--17983
"111110001000001001110011100000000000",--17984
"001111000100000010000000000000000010",--17985
"111110001010001010000100000000000000",--17986
"001101000010000000100000000000000011",--17987
"011100000101000000000000000000000100",--17988
"001011000000000001100000000100100110",--17989
"001011000000000001110000000100100111",--17990
"001011000000000010000000000100101000",--17991
"000101000000000000000100011001100101",--17992
"001101000010000000100000000000001001",--17993
"001111000100000010010000000000000010",--17994
"111110001000001010010100100000000000",--17995
"001111000100000010100000000000000001",--17996
"111110001010001010100101000000000000",--17997
"111110010010000010100100100000000000",--17998
"101111000001110010100011111100000000",--17999
"111110010010001010100100100000000000",--18000
"111110001100000010010011000000000000",--18001
"001011000000000001100000000100100110",--18002
"001111000100000001100000000000000010",--18003
"111110000110001001100011000000000000",--18004
"001111000100000010010000000000000000",--18005
"111110001010001010010010100000000000",--18006
"111110001100000001010010100000000000",--18007
"101111000001110001100011111100000000",--18008
"111110001010001001100010100000000000",--18009
"111110001110000001010010100000000000",--18010
"001011000000000001010000000100100111",--18011
"001111000100000001010000000000000001",--18012
"111110000110001001010001100000000000",--18013
"001111000100000001010000000000000000",--18014
"111110001000001001010010000000000000",--18015
"111110000110000001000001100000000000",--18016
"101111000001110001000011111100000000",--18017
"111110000110001001000001100000000000",--18018
"111110010000000000110001100000000000",--18019
"001011000000000000110000000100101000",--18020
"001111000000000000110000000100100110",--18021
"111110000110001000110001100000000000",--18022
"001111000000000001000000000100100111",--18023
"111110001000001001000010000000000000",--18024
"111110000110000001000001100000000000",--18025
"001111000000000001000000000100101000",--18026
"111110001000001001000010000000000000",--18027
"111110000110000001000001100000000000",--18028
"111110000110100000000001100000000000",--18029
"011110000111000000000000000000000010",--18030
"101110000011111000000001100000000000",--18031
"000101000000000000000100011001110110",--18032
"001101000010000000100000000000000110",--18033
"011100000101000000000000000000000010",--18034
"111110000110011000000001100000000000",--18035
"000101000000000000000100011001110110",--18036
"111110000110011000000001100000000010",--18037
"001111000000000001000000000100100110",--18038
"111110001000001000110010000000000000",--18039
"001011000000000001000000000100100110",--18040
"001111000000000001000000000100100111",--18041
"111110001000001000110010000000000000",--18042
"001011000000000001000000000100100111",--18043
"001111000000000001000000000100101000",--18044
"111110001000001000110001100000000000",--18045
"001011000000000000110000000100101000",--18046
"001101000010000000100000000000000000",--18047
"001101000010000000110000000000001000",--18048
"001111000110000000110000000000000000",--18049
"001011000000000000110000000100100011",--18050
"001111000110000000110000000000000001",--18051
"001011000000000000110000000100100100",--18052
"001111000110000000110000000000000010",--18053
"001011000000000000110000000100100101",--18054
"001001111100000000011111111111111000",--18055
"011111000101000000010000000000100011",--18056
"001111000000000000110000000100101010",--18057
"001101000010000000100000000000000101",--18058
"001111000100000001000000000000000000",--18059
"111110000110010001000001100000000000",--18060
"101111001001110001000011110101001100",--18061
"101111001001100001001100110011001101",--18062
"111110000110001001000010000000000000",--18063
"101110001000110000000010000000000000",--18064
"101111000001110001010100000110100000",--18065
"111110001000001001010010000000000000",--18066
"111110000110010001000001100000000000",--18067
"101111000001110001000100000100100000",--18068
"001111000000000001010000000100101100",--18069
"001111000100000001100000000000000010",--18070
"111110001010010001100010100000000000",--18071
"101111001101110001100011110101001100",--18072
"101111001101100001101100110011001101",--18073
"111110001010001001100011000000000000",--18074
"101110001100110000000011000000000000",--18075
"101111000001110001110100000110100000",--18076
"111110001100001001110011000000000000",--18077
"111110001010010001100010100000000000",--18078
"101111000001110001100100000100100000",--18079
"010110001001000000110000000000000101",--18080
"010110001101000001010000000000000010",--18081
"101111000001110000110100001101111111",--18082
"000101000000000000000100011010101010",--18083
"101110000001111000000001100000000000",--18084
"000101000000000000000100011010101010",--18085
"010110001101000001010000000000000010",--18086
"101110000001111000000001100000000000",--18087
"000101000000000000000100011010101010",--18088
"101111000001110000110100001101111111",--18089
"001011000000000000110000000100100100",--18090
"000101000000000000000100011111100101",--18091
"011111000101000000100000000000001111",--18092
"001111000000000000110000000100101011",--18093
"101111000001110001000011111010000000",--18094
"111110000110001001000001100000000000",--18095
"001001111100000111111111111111110111",--18096
"000111000000000000000111011000000010",--18097
"001101111100000111111111111111110111",--18098
"111110000110001000110001100000000000",--18099
"101111000001110001000100001101111111",--18100
"111110001000001000110010000000000000",--18101
"001011000000000001000000000100100011",--18102
"101111000001110001000100001101111111",--18103
"111110000110010000010001100000000010",--18104
"111110001000001000110001100000000000",--18105
"001011000000000000110000000100100100",--18106
"000101000000000000000100011111100101",--18107
"011111000101000000110000000000011111",--18108
"001111000000000000110000000100101010",--18109
"001101000010000000100000000000000101",--18110
"001111000100000001000000000000000000",--18111
"111110000110010001000001100000000000",--18112
"001111000000000001000000000100101100",--18113
"001111000100000001010000000000000010",--18114
"111110001000010001010010000000000000",--18115
"111110000110001000110001100000000000",--18116
"111110001000001001000010000000000000",--18117
"111110000110000001000001100000000000",--18118
"111110000110100000000001100000000000",--18119
"101111001001110001000011110111001100",--18120
"101111001001100001001100110011001100",--18121
"111110000110001001000001100000000000",--18122
"101110000110110000000010000000000000",--18123
"111110000110010001000001100000000000",--18124
"101111001001110001000100000001001001",--18125
"101111001001100001000000111111011011",--18126
"111110000110001001000001100000000000",--18127
"001001111100000111111111111111110111",--18128
"000111000000000000000111010110111000",--18129
"001101111100000111111111111111110111",--18130
"111110000110001000110001100000000000",--18131
"101111000001110001000100001101111111",--18132
"111110000110001001000010000000000000",--18133
"001011000000000001000000000100100100",--18134
"111110000110010000010001100000000010",--18135
"101111000001110001000100001101111111",--18136
"111110000110001001000001100000000000",--18137
"001011000000000000110000000100100101",--18138
"000101000000000000000100011111100101",--18139
"011111000101000001000000000100001000",--18140
"001111000000000000110000000100101010",--18141
"001101000010000000100000000000000101",--18142
"001111000100000001000000000000000000",--18143
"111110000110010001000001100000000000",--18144
"001101000010000000110000000000000100",--18145
"001111000110000001000000000000000000",--18146
"111110001000100000000010000000000000",--18147
"111110000110001001000001100000000000",--18148
"001111000000000001000000000100101100",--18149
"001111000100000001010000000000000010",--18150
"111110001000010001010010000000000000",--18151
"001111000110000001010000000000000010",--18152
"111110001010100000000010100000000000",--18153
"111110001000001001010010000000000000",--18154
"111110000110001000110010100000000000",--18155
"111110001000001001000011000000000000",--18156
"111110001010000001100010100000000000",--18157
"101110000111111000000011000000000001",--18158
"101111001111110001110011100011010001",--18159
"101111001111100001111011011100010111",--18160
"001001111100000000111111111111110111",--18161
"001001111100000000101111111111110110",--18162
"001011111100000001011111111111110101",--18163
"010110001111000001100000000000000010",--18164
"101111000001110000110100000101110000",--18165
"000101000000000000000100011101011010",--18166
"111110000110011000000001100000000000",--18167
"111110001000001000110001100000000001",--18168
"010110000111000000010000000000000010",--18169
"101001000000000001000000000000000001",--18170
"000101000000000000000100011100000001",--18171
"011010000111000000100000000000000010",--18172
"101001000000000001001111111111111111",--18173
"000101000000000000000100011100000001",--18174
"101000000001111000000010000000000000",--18175
"000101000000000000000100011100000010",--18176
"111110000110011000000001100000000000",--18177
"111110000110001000110010000000000000",--18178
"101111000001110001100100001011110010",--18179
"111110001100001001000011000000000000",--18180
"101111001111110001110011110100110010",--18181
"101111001111100001110001011001000011",--18182
"111110001100001001110011000000000000",--18183
"101111000001110001110100001011001000",--18184
"111110001110001001000011100000000000",--18185
"101111000001110010000100000110101000",--18186
"111110010000000001100011000000000000",--18187
"111110001100011000000011000000000000",--18188
"111110001110001001100011000000000000",--18189
"101111000001110001110100001010100010",--18190
"111110001110001001000011100000000000",--18191
"101111000001110010000100000110011000",--18192
"111110010000000001100011000000000000",--18193
"111110001100011000000011000000000000",--18194
"111110001110001001100011000000000000",--18195
"101111000001110001110100001010000000",--18196
"111110001110001001000011100000000000",--18197
"101111000001110010000100000110001000",--18198
"111110010000000001100011000000000000",--18199
"111110001100011000000011000000000000",--18200
"111110001110001001100011000000000000",--18201
"101111000001110001110100001001000100",--18202
"111110001110001001000011100000000000",--18203
"101111000001110010000100000101110000",--18204
"111110010000000001100011000000000000",--18205
"111110001100011000000011000000000000",--18206
"111110001110001001100011000000000000",--18207
"101111000001110001110100001000010000",--18208
"111110001110001001000011100000000000",--18209
"101111000001110010000100000101010000",--18210
"111110010000000001100011000000000000",--18211
"111110001100011000000011000000000000",--18212
"111110001110001001100011000000000000",--18213
"101111000001110001110100000111001000",--18214
"111110001110001001000011100000000000",--18215
"101111000001110010000100000100110000",--18216
"111110010000000001100011000000000000",--18217
"111110001100011000000011000000000000",--18218
"111110001110001001100011000000000000",--18219
"101111000001110001110100000110000000",--18220
"111110001110001001000011100000000000",--18221
"101111000001110010000100000100010000",--18222
"111110010000000001100011000000000000",--18223
"111110001100011000000011000000000000",--18224
"111110001110001001100011000000000000",--18225
"101111000001110001110100000100010000",--18226
"111110001110001001000011100000000000",--18227
"101111000001110010000100000011100000",--18228
"111110010000000001100011000000000000",--18229
"111110001100011000000011000000000000",--18230
"111110001110001001100011000000000000",--18231
"101111000001110010000100000010000000",--18232
"111110010000001001000100000000000000",--18233
"101111000001110010010100000010100000",--18234
"111110010010000001100011000000000000",--18235
"111110001100011000000011000000000000",--18236
"111110010000001001100011000000000000",--18237
"001001111100000001001111111111110100",--18238
"001011111100000000111111111111110011",--18239
"101110001101111000000010100000000000",--18240
"101110000011111000000001100000000000",--18241
"001001111100000111111111111111110010",--18242
"101001111100010111100000000000001111",--18243
"000111000000000000000000001101001100",--18244
"101001111100000111100000000000001111",--18245
"001101111100000111111111111111110010",--18246
"111110000110000000010001100000000000",--18247
"111110000110011000000001100000000000",--18248
"001111111100000001001111111111110011",--18249
"111110001000001000110001100000000000",--18250
"001101111100000000011111111111110100",--18251
"010100000011000000000000000000000100",--18252
"101111001001110001000011111111001001",--18253
"101111001001100001000000111111011010",--18254
"111110001000010000110001100000000000",--18255
"000101000000000000000100011101010101",--18256
"011000000011000000000000000000000011",--18257
"101111001001110001001011111111001001",--18258
"101111001001100001000000111111011010",--18259
"111110001000010000110001100000000000",--18260
"101111000001110001000100000111110000",--18261
"111110000110001001000001100000000000",--18262
"101111001001110001000011111010100010",--18263
"101111001001100001001111100110000010",--18264
"111110000110001001000001100000000000",--18265
"101110000110110000000010000000000000",--18266
"111110000110010001000001100000000000",--18267
"001111111100000001001111111111110101",--18268
"101110001001111000000010100000000001",--18269
"101111001101110001100011100011010001",--18270
"101111001101100001101011011100010111",--18271
"001011111100000000111111111111110100",--18272
"010110001101000001010000000000000010",--18273
"101111000001110000110100000101110000",--18274
"000101000000000000000100011111010000",--18275
"001111000000000001010000000100101011",--18276
"001101111100000000011111111111110110",--18277
"001111000010000001100000000000000001",--18278
"111110001010010001100010100000000000",--18279
"001101111100000000011111111111110111",--18280
"001111000010000001100000000000000001",--18281
"111110001100100000000011000000000000",--18282
"111110001010001001100010100000000000",--18283
"111110001000011000000010000000000000",--18284
"111110001010001001000010000000000001",--18285
"010110001001000000010000000000000010",--18286
"101001000000000000010000000000000001",--18287
"000101000000000000000100011101110110",--18288
"011010001001000000100000000000000010",--18289
"101001000000000000011111111111111111",--18290
"000101000000000000000100011101110110",--18291
"101000000001111000000000100000000000",--18292
"000101000000000000000100011101110111",--18293
"111110001000011000000010000000000000",--18294
"111110001000001001000010100000000000",--18295
"101111000001110001100100001011110010",--18296
"111110001100001001010011000000000000",--18297
"101111001111110001110011110100110010",--18298
"101111001111100001110001011001000011",--18299
"111110001100001001110011000000000000",--18300
"101111000001110001110100001011001000",--18301
"111110001110001001010011100000000000",--18302
"101111000001110010000100000110101000",--18303
"111110010000000001100011000000000000",--18304
"111110001100011000000011000000000000",--18305
"111110001110001001100011000000000000",--18306
"101111000001110001110100001010100010",--18307
"111110001110001001010011100000000000",--18308
"101111000001110010000100000110011000",--18309
"111110010000000001100011000000000000",--18310
"111110001100011000000011000000000000",--18311
"111110001110001001100011000000000000",--18312
"101111000001110001110100001010000000",--18313
"111110001110001001010011100000000000",--18314
"101111000001110010000100000110001000",--18315
"111110010000000001100011000000000000",--18316
"111110001100011000000011000000000000",--18317
"111110001110001001100011000000000000",--18318
"101111000001110001110100001001000100",--18319
"111110001110001001010011100000000000",--18320
"101111000001110010000100000101110000",--18321
"111110010000000001100011000000000000",--18322
"111110001100011000000011000000000000",--18323
"111110001110001001100011000000000000",--18324
"101111000001110001110100001000010000",--18325
"111110001110001001010011100000000000",--18326
"101111000001110010000100000101010000",--18327
"111110010000000001100011000000000000",--18328
"111110001100011000000011000000000000",--18329
"111110001110001001100011000000000000",--18330
"101111000001110001110100000111001000",--18331
"111110001110001001010011100000000000",--18332
"101111000001110010000100000100110000",--18333
"111110010000000001100011000000000000",--18334
"111110001100011000000011000000000000",--18335
"111110001110001001100011000000000000",--18336
"101111000001110001110100000110000000",--18337
"111110001110001001010011100000000000",--18338
"101111000001110010000100000100010000",--18339
"111110010000000001100011000000000000",--18340
"111110001100011000000011000000000000",--18341
"111110001110001001100011000000000000",--18342
"101111000001110001110100000100010000",--18343
"111110001110001001010011100000000000",--18344
"101111000001110010000100000011100000",--18345
"111110010000000001100011000000000000",--18346
"111110001100011000000011000000000000",--18347
"111110001110001001100011000000000000",--18348
"101111000001110010000100000010000000",--18349
"111110010000001001010100000000000000",--18350
"101111000001110010010100000010100000",--18351
"111110010010000001100011000000000000",--18352
"111110001100011000000011000000000000",--18353
"111110010000001001100011000000000000",--18354
"001001111100000000011111111111110011",--18355
"001011111100000001001111111111110010",--18356
"101110001011111000000010000000000000",--18357
"101110000011111000000001100000000000",--18358
"101110001101111000000010100000000000",--18359
"001001111100000111111111111111110001",--18360
"101001111100010111100000000000010000",--18361
"000111000000000000000000001101001100",--18362
"101001111100000111100000000000010000",--18363
"001101111100000111111111111111110001",--18364
"111110000110000000010001100000000000",--18365
"111110000110011000000001100000000000",--18366
"001111111100000001001111111111110010",--18367
"111110001000001000110001100000000000",--18368
"001101111100000000011111111111110011",--18369
"010100000011000000000000000000000100",--18370
"101111001001110001000011111111001001",--18371
"101111001001100001000000111111011010",--18372
"111110001000010000110001100000000000",--18373
"000101000000000000000100011111001011",--18374
"011000000011000000000000000000000011",--18375
"101111001001110001001011111111001001",--18376
"101111001001100001000000111111011010",--18377
"111110001000010000110001100000000000",--18378
"101111000001110001000100000111110000",--18379
"111110000110001001000001100000000000",--18380
"101111001001110001000011111010100010",--18381
"101111001001100001001111100110000010",--18382
"111110000110001001000001100000000000",--18383
"101110000110110000000010000000000000",--18384
"111110000110010001000001100000000000",--18385
"101111001001110001000011111000011001",--18386
"101111001001100001001001100110011010",--18387
"101111000001110001010011111100000000",--18388
"001111111100000001101111111111110100",--18389
"111110001010010001100010100000000000",--18390
"111110001010001001010010100000000000",--18391
"111110001000010001010010000000000000",--18392
"101111000001110001010011111100000000",--18393
"111110001010010000110001100000000000",--18394
"111110000110001000110001100000000000",--18395
"111110001000010000110001100000000000",--18396
"011010000111000000000000000000000001",--18397
"101110000001111000000001100000000000",--18398
"101111000001110001000100001101111111",--18399
"111110001000001000110001100000000000",--18400
"101111001001110001000100000001010101",--18401
"101111001001100001000101010101010101",--18402
"111110000110001001000001100000000000",--18403
"001011000000000000110000000100100101",--18404
"001101000000000000100000000100110000",--18405
"001101000100000000010000000000000000",--18406
"001101000010000000110000000000000000",--18407
"010011000111000000000000000010110100",--18408
"001001111100000000011111111111110111",--18409
"001001111100000000101111111111110110",--18410
"010011000111011000110000000010100010",--18411
"001101000110000001000000000101101101",--18412
"001111000000000000110000000100101010",--18413
"001101001000000001010000000000000101",--18414
"001111001010000001000000000000000000",--18415
"111110000110010001000001100000000000",--18416
"001111000000000001000000000100101011",--18417
"001111001010000001010000000000000001",--18418
"111110001000010001010010000000000000",--18419
"001111000000000001010000000100101100",--18420
"001111001010000001100000000000000010",--18421
"111110001010010001100010100000000000",--18422
"001101000110000000110000000010111110",--18423
"001101001000000001010000000000000001",--18424
"011111001011000000010000000000110111",--18425
"001111000110000001100000000000000000",--18426
"111110001100010000110011000000000000",--18427
"001111000110000001110000000000000001",--18428
"111110001100001001110011000000000000",--18429
"001111000000000001110000000011111011",--18430
"111110001100001001110011100000000000",--18431
"111110001110000001000011100000000001",--18432
"001101001000000001000000000000000100",--18433
"001111001000000010000000000000000001",--18434
"010110010001000001110000000000000111",--18435
"001111000000000001110000000011111100",--18436
"111110001100001001110011100000000000",--18437
"111110001110000001010011100000000001",--18438
"001111001000000010000000000000000010",--18439
"010110010001000001110000000000000010",--18440
"001111000110000001110000000000000001",--18441
"011110001111000000000000000000100100",--18442
"001111000110000001100000000000000010",--18443
"111110001100010001000011000000000000",--18444
"001111000110000001110000000000000011",--18445
"111110001100001001110011000000000000",--18446
"001111000000000001110000000011111010",--18447
"111110001100001001110011100000000000",--18448
"111110001110000000110011100000000001",--18449
"001111001000000010000000000000000000",--18450
"010110010001000001110000000000000111",--18451
"001111000000000001110000000011111100",--18452
"111110001100001001110011100000000000",--18453
"111110001110000001010011100000000001",--18454
"001111001000000010000000000000000010",--18455
"010110010001000001110000000000000010",--18456
"001111000110000001110000000000000011",--18457
"011110001111000000000000000000010010",--18458
"001111000110000001100000000000000100",--18459
"111110001100010001010010100000000000",--18460
"001111000110000001100000000000000101",--18461
"111110001010001001100010100000000000",--18462
"001111000000000001100000000011111010",--18463
"111110001010001001100011000000000000",--18464
"111110001100000000110001100000000001",--18465
"001111001000000001100000000000000000",--18466
"010110001101000000110000000001100001",--18467
"001111000000000000110000000011111011",--18468
"111110001010001000110001100000000000",--18469
"111110000110000001000001100000000001",--18470
"001111001000000001000000000000000001",--18471
"010110001001000000110000000001011100",--18472
"001111000110000000110000000000000101",--18473
"010010000111000000000000000001011010",--18474
"001011000000000001010000000100101111",--18475
"000101000000000000000100100001111001",--18476
"001011000000000001100000000100101111",--18477
"000101000000000000000100100001111001",--18478
"001011000000000001100000000100101111",--18479
"000101000000000000000100100001111001",--18480
"011111001011000000100000000000001100",--18481
"001111000110000001100000000000000000",--18482
"011010001101000000000000000001010001",--18483
"001111000110000001100000000000000001",--18484
"111110001100001000110001100000000000",--18485
"001111000110000001100000000000000010",--18486
"111110001100001001000010000000000000",--18487
"111110000110000001000001100000000000",--18488
"001111000110000001000000000000000011",--18489
"111110001000001001010010000000000000",--18490
"111110000110000001000001100000000000",--18491
"001011000000000000110000000100101111",--18492
"000101000000000000000100100001111001",--18493
"001111000110000001100000000000000000",--18494
"010010001101000000000000000001000101",--18495
"001111000110000001110000000000000001",--18496
"111110001110001000110011100000000000",--18497
"001111000110000010000000000000000010",--18498
"111110010000001001000100000000000000",--18499
"111110001110000010000011100000000000",--18500
"001111000110000010000000000000000011",--18501
"111110010000001001010100000000000000",--18502
"111110001110000010000011100000000000",--18503
"111110000110001000110100000000000000",--18504
"001101001000000001100000000000000100",--18505
"001111001100000010010000000000000000",--18506
"111110010000001010010100000000000000",--18507
"111110001000001001000100100000000000",--18508
"001111001100000010100000000000000001",--18509
"111110010010001010100100100000000000",--18510
"111110010000000010010100000000000000",--18511
"111110001010001001010100100000000000",--18512
"001111001100000010100000000000000010",--18513
"111110010010001010100100100000000000",--18514
"111110010000000010010100000000000000",--18515
"001101001000000001100000000000000011",--18516
"011100001101000000000000000000000011",--18517
"101110010001111000000001100000000000",--18518
"011111001011000000110000000000010000",--18519
"000101000000000000000100100001100111",--18520
"111110001000001001010100100000000000",--18521
"001101001000000001100000000000001001",--18522
"001111001100000010100000000000000000",--18523
"111110010010001010100100100000000000",--18524
"111110010000000010010100000000000000",--18525
"111110001010001000110010100000000000",--18526
"001111001100000010010000000000000001",--18527
"111110001010001010010010100000000000",--18528
"111110010000000001010010100000000000",--18529
"111110000110001001000001100000000000",--18530
"001111001100000001000000000000000010",--18531
"111110000110001001000001100000000000",--18532
"111110001010000000110001100000000000",--18533
"011111001011000000110000000000000001",--18534
"111110000110010000010001100000000000",--18535
"111110001110001001110010000000000000",--18536
"111110001100001000110001100000000000",--18537
"111110001000010000110001100000000000",--18538
"010110000111000000000000000000011001",--18539
"001101001000000001000000000000000110",--18540
"011100001001000000000000000000000110",--18541
"111110000110100000000001100000000000",--18542
"111110001110010000110001100000000000",--18543
"001111000110000001000000000000000100",--18544
"111110000110001001000001100000000000",--18545
"001011000000000000110000000100101111",--18546
"000101000000000000000100100001111001",--18547
"111110000110100000000001100000000000",--18548
"111110001110000000110001100000000000",--18549
"001111000110000001000000000000000100",--18550
"111110000110001001000001100000000000",--18551
"001011000000000000110000000100101111",--18552
"001111000000000000110000000100101111",--18553
"101111001001110001001011110111001100",--18554
"101111001001100001001100110011001101",--18555
"010110001001000000110000000000001000",--18556
"101000000011111000000001000000000000",--18557
"101001000000000000010000000000000001",--18558
"001001111100000111111111111111110101",--18559
"101001111100010111100000000000001100",--18560
"000111000000000000000000110101111110",--18561
"101001111100000111100000000000001100",--18562
"001101111100000111111111111111110101",--18563
"011100000011000000000000000000001001",--18564
"101001000000000000010000000000000001",--18565
"001101111100000000101111111111110110",--18566
"001001111100000111111111111111110101",--18567
"101001111100010111100000000000001100",--18568
"000111000000000000000000111111111011",--18569
"101001111100000111100000000000001100",--18570
"001101111100000111111111111111110101",--18571
"011100000011000000000000001011111100",--18572
"000101000000000000000100100010011101",--18573
"101001000000000000010000000000000001",--18574
"001101111100000000101111111111110111",--18575
"001001111100000111111111111111110101",--18576
"101001111100010111100000000000001100",--18577
"000111000000000000000000110101111110",--18578
"101001111100000111100000000000001100",--18579
"001101111100000111111111111111110101",--18580
"011100000011000000000000001011110011",--18581
"101001000000000000010000000000000001",--18582
"001101111100000000101111111111110110",--18583
"101001111100010111100000000000001100",--18584
"000111000000000000000000111111111011",--18585
"101001111100000111100000000000001100",--18586
"001101111100000111111111111111110101",--18587
"011100000011000000000000001011101100",--18588
"101111000111110000111011101111011010",--18589
"101111000111100000110111010000001101",--18590
"001111111100000001001111111111111010",--18591
"111110001000001000110001100000000000",--18592
"001111000000000001000000000100100110",--18593
"001111000000000001010000000101100100",--18594
"111110001000001001010010000000000000",--18595
"001111000000000001010000000100100111",--18596
"001111000000000001100000000101100101",--18597
"111110001010001001100010100000000000",--18598
"111110001000000001010010000000000000",--18599
"001111000000000001010000000100101000",--18600
"001111000000000001100000000101100110",--18601
"111110001010001001100010100000000000",--18602
"111110001000000001010010000000000010",--18603
"010110001001000000000000000000000001",--18604
"000101000000000000000100100010101111",--18605
"101110000001111000000010000000000000",--18606
"111110000110001001000001100000000000",--18607
"001101111100000000011111111111111000",--18608
"001101000010000000010000000000000111",--18609
"001111000010000001000000000000000000",--18610
"111110000110001001000001100000000000",--18611
"001111000000000001000000000100100000",--18612
"001111000000000001010000000100100011",--18613
"111110000110001001010010100000000000",--18614
"111110001000000001010010000000000000",--18615
"001011000000000001000000000100100000",--18616
"001111000000000001000000000100100001",--18617
"001111000000000001010000000100100100",--18618
"111110000110001001010010100000000000",--18619
"111110001000000001010010000000000000",--18620
"001011000000000001000000000100100001",--18621
"001111000000000001000000000100100010",--18622
"001111000000000001010000000100100101",--18623
"111110000110001001010001100000000000",--18624
"111110001000000000110001100000000000",--18625
"001011000000000000110000000100100010",--18626
"000101000000000000000100101110001001",--18627
"001100000110000000010001100000000000",--18628
"101111001001110001000100111001101110",--18629
"101111001001100001000110101100101000",--18630
"001011000000000001000000000100101101",--18631
"001101000000000000100000000100110000",--18632
"001011111100000000111111111111111010",--18633
"001001111100000000111111111111111001",--18634
"101000000001111000000000100000000000",--18635
"001001111100000111111111111111111000",--18636
"101001111100010111100000000000001001",--18637
"000111000000000000000010110111111111",--18638
"101001111100000111100000000000001001",--18639
"001101111100000111111111111111111000",--18640
"001111000000000000110000000100101101",--18641
"101111001001110001001011110111001100",--18642
"101111001001100001001100110011001101",--18643
"010110000111000001000000001010110100",--18644
"101111001001110001000100110010111110",--18645
"101111001001100001001011110000100000",--18646
"010110001001000000110000001010110001",--18647
"001101000000000000010000000100101001",--18648
"001101000010000000010000000101101101",--18649
"001101000010000000100000000000000001",--18650
"011111000101000000010000000000010011",--18651
"001101111100000000101111111111111001",--18652
"001101000100000000100000000000000000",--18653
"001101000000000000110000000100101110",--18654
"001011000000000000000000000100100110",--18655
"001011000000000000000000000100100111",--18656
"001011000000000000000000000100101000",--18657
"101001000110010001000000000000000001",--18658
"101001000110010000110000000000000001",--18659
"001110000100000000110001100000000000",--18660
"011110000111000000000000000000000010",--18661
"101110000001111000000001100000000000",--18662
"000101000000000000000100100011101100",--18663
"010110000111000000000000000000000010",--18664
"101110000011111000000001100000000000",--18665
"000101000000000000000100100011101100",--18666
"101110000101111000000001100000000000",--18667
"101110000111111000000001100000000010",--18668
"001011001000000000110000000100100110",--18669
"000101000000000000000100100101000101",--18670
"011111000101000000100000000000001000",--18671
"001101000010000000100000000000000100",--18672
"001111000100010000110000000000000000",--18673
"001011000000000000110000000100100110",--18674
"001111000100010000110000000000000001",--18675
"001011000000000000110000000100100111",--18676
"001111000100010000110000000000000010",--18677
"001011000000000000110000000100101000",--18678
"000101000000000000000100100101000101",--18679
"001111000000000000110000000100101010",--18680
"001101000010000000100000000000000101",--18681
"001111000100000001000000000000000000",--18682
"111110000110010001000001100000000000",--18683
"001111000000000001000000000100101011",--18684
"001111000100000001010000000000000001",--18685
"111110001000010001010010000000000000",--18686
"001111000000000001010000000100101100",--18687
"001111000100000001100000000000000010",--18688
"111110001010010001100010100000000000",--18689
"001101000010000000100000000000000100",--18690
"001111000100000001100000000000000000",--18691
"111110000110001001100011000000000000",--18692
"001111000100000001110000000000000001",--18693
"111110001000001001110011100000000000",--18694
"001111000100000010000000000000000010",--18695
"111110001010001010000100000000000000",--18696
"001101000010000000100000000000000011",--18697
"011100000101000000000000000000000100",--18698
"001011000000000001100000000100100110",--18699
"001011000000000001110000000100100111",--18700
"001011000000000010000000000100101000",--18701
"000101000000000000000100100100101011",--18702
"001101000010000000100000000000001001",--18703
"001111000100000010010000000000000010",--18704
"111110001000001010010100100000000000",--18705
"001111000100000010100000000000000001",--18706
"111110001010001010100101000000000000",--18707
"111110010010000010100100100000000000",--18708
"101111000001110010100011111100000000",--18709
"111110010010001010100100100000000000",--18710
"111110001100000010010011000000000000",--18711
"001011000000000001100000000100100110",--18712
"001111000100000001100000000000000010",--18713
"111110000110001001100011000000000000",--18714
"001111000100000010010000000000000000",--18715
"111110001010001010010010100000000000",--18716
"111110001100000001010010100000000000",--18717
"101111000001110001100011111100000000",--18718
"111110001010001001100010100000000000",--18719
"111110001110000001010010100000000000",--18720
"001011000000000001010000000100100111",--18721
"001111000100000001010000000000000001",--18722
"111110000110001001010001100000000000",--18723
"001111000100000001010000000000000000",--18724
"111110001000001001010010000000000000",--18725
"111110000110000001000001100000000000",--18726
"101111000001110001000011111100000000",--18727
"111110000110001001000001100000000000",--18728
"111110010000000000110001100000000000",--18729
"001011000000000000110000000100101000",--18730
"001111000000000000110000000100100110",--18731
"111110000110001000110001100000000000",--18732
"001111000000000001000000000100100111",--18733
"111110001000001001000010000000000000",--18734
"111110000110000001000001100000000000",--18735
"001111000000000001000000000100101000",--18736
"111110001000001001000010000000000000",--18737
"111110000110000001000001100000000000",--18738
"111110000110100000000001100000000000",--18739
"011110000111000000000000000000000010",--18740
"101110000011111000000001100000000000",--18741
"000101000000000000000100100100111100",--18742
"001101000010000000100000000000000110",--18743
"011100000101000000000000000000000010",--18744
"111110000110011000000001100000000000",--18745
"000101000000000000000100100100111100",--18746
"111110000110011000000001100000000010",--18747
"001111000000000001000000000100100110",--18748
"111110001000001000110010000000000000",--18749
"001011000000000001000000000100100110",--18750
"001111000000000001000000000100100111",--18751
"111110001000001000110010000000000000",--18752
"001011000000000001000000000100100111",--18753
"001111000000000001000000000100101000",--18754
"111110001000001000110001100000000000",--18755
"001011000000000000110000000100101000",--18756
"001101000010000000100000000000000000",--18757
"001101000010000000110000000000001000",--18758
"001111000110000000110000000000000000",--18759
"001011000000000000110000000100100011",--18760
"001111000110000000110000000000000001",--18761
"001011000000000000110000000100100100",--18762
"001111000110000000110000000000000010",--18763
"001011000000000000110000000100100101",--18764
"001001111100000000011111111111111000",--18765
"011111000101000000010000000000100011",--18766
"001111000000000000110000000100101010",--18767
"001101000010000000100000000000000101",--18768
"001111000100000001000000000000000000",--18769
"111110000110010001000001100000000000",--18770
"101111001001110001000011110101001100",--18771
"101111001001100001001100110011001101",--18772
"111110000110001001000010000000000000",--18773
"101110001000110000000010000000000000",--18774
"101111000001110001010100000110100000",--18775
"111110001000001001010010000000000000",--18776
"111110000110010001000001100000000000",--18777
"101111000001110001000100000100100000",--18778
"001111000000000001010000000100101100",--18779
"001111000100000001100000000000000010",--18780
"111110001010010001100010100000000000",--18781
"101111001101110001100011110101001100",--18782
"101111001101100001101100110011001101",--18783
"111110001010001001100011000000000000",--18784
"101110001100110000000011000000000000",--18785
"101111000001110001110100000110100000",--18786
"111110001100001001110011000000000000",--18787
"111110001010010001100010100000000000",--18788
"101111000001110001100100000100100000",--18789
"010110001001000000110000000000000101",--18790
"010110001101000001010000000000000010",--18791
"101111000001110000110100001101111111",--18792
"000101000000000000000100100101110000",--18793
"101110000001111000000001100000000000",--18794
"000101000000000000000100100101110000",--18795
"010110001101000001010000000000000010",--18796
"101110000001111000000001100000000000",--18797
"000101000000000000000100100101110000",--18798
"101111000001110000110100001101111111",--18799
"001011000000000000110000000100100100",--18800
"000101000000000000000100101010101011",--18801
"011111000101000000100000000000001111",--18802
"001111000000000000110000000100101011",--18803
"101111000001110001000011111010000000",--18804
"111110000110001001000001100000000000",--18805
"001001111100000111111111111111110111",--18806
"000111000000000000000111011000000010",--18807
"001101111100000111111111111111110111",--18808
"111110000110001000110001100000000000",--18809
"101111000001110001000100001101111111",--18810
"111110001000001000110010000000000000",--18811
"001011000000000001000000000100100011",--18812
"101111000001110001000100001101111111",--18813
"111110000110010000010001100000000010",--18814
"111110001000001000110001100000000000",--18815
"001011000000000000110000000100100100",--18816
"000101000000000000000100101010101011",--18817
"011111000101000000110000000000011111",--18818
"001111000000000000110000000100101010",--18819
"001101000010000000100000000000000101",--18820
"001111000100000001000000000000000000",--18821
"111110000110010001000001100000000000",--18822
"001111000000000001000000000100101100",--18823
"001111000100000001010000000000000010",--18824
"111110001000010001010010000000000000",--18825
"111110000110001000110001100000000000",--18826
"111110001000001001000010000000000000",--18827
"111110000110000001000001100000000000",--18828
"111110000110100000000001100000000000",--18829
"101111001001110001000011110111001100",--18830
"101111001001100001001100110011001100",--18831
"111110000110001001000001100000000000",--18832
"101110000110110000000010000000000000",--18833
"111110000110010001000001100000000000",--18834
"101111001001110001000100000001001001",--18835
"101111001001100001000000111111011011",--18836
"111110000110001001000001100000000000",--18837
"001001111100000111111111111111110111",--18838
"000111000000000000000111010110111000",--18839
"001101111100000111111111111111110111",--18840
"111110000110001000110001100000000000",--18841
"101111000001110001000100001101111111",--18842
"111110000110001001000010000000000000",--18843
"001011000000000001000000000100100100",--18844
"111110000110010000010001100000000010",--18845
"101111000001110001000100001101111111",--18846
"111110000110001001000001100000000000",--18847
"001011000000000000110000000100100101",--18848
"000101000000000000000100101010101011",--18849
"011111000101000001000000000100001000",--18850
"001111000000000000110000000100101010",--18851
"001101000010000000100000000000000101",--18852
"001111000100000001000000000000000000",--18853
"111110000110010001000001100000000000",--18854
"001101000010000000110000000000000100",--18855
"001111000110000001000000000000000000",--18856
"111110001000100000000010000000000000",--18857
"111110000110001001000001100000000000",--18858
"001111000000000001000000000100101100",--18859
"001111000100000001010000000000000010",--18860
"111110001000010001010010000000000000",--18861
"001111000110000001010000000000000010",--18862
"111110001010100000000010100000000000",--18863
"111110001000001001010010000000000000",--18864
"111110000110001000110010100000000000",--18865
"111110001000001001000011000000000000",--18866
"111110001010000001100010100000000000",--18867
"101110000111111000000011000000000001",--18868
"101111001111110001110011100011010001",--18869
"101111001111100001111011011100010111",--18870
"001001111100000000111111111111110111",--18871
"001001111100000000101111111111110110",--18872
"001011111100000001011111111111110101",--18873
"010110001111000001100000000000000010",--18874
"101111000001110000110100000101110000",--18875
"000101000000000000000100101000100000",--18876
"111110000110011000000001100000000000",--18877
"111110001000001000110001100000000001",--18878
"010110000111000000010000000000000010",--18879
"101001000000000001000000000000000001",--18880
"000101000000000000000100100111000111",--18881
"011010000111000000100000000000000010",--18882
"101001000000000001001111111111111111",--18883
"000101000000000000000100100111000111",--18884
"101000000001111000000010000000000000",--18885
"000101000000000000000100100111001000",--18886
"111110000110011000000001100000000000",--18887
"111110000110001000110010000000000000",--18888
"101111000001110001100100001011110010",--18889
"111110001100001001000011000000000000",--18890
"101111001111110001110011110100110010",--18891
"101111001111100001110001011001000011",--18892
"111110001100001001110011000000000000",--18893
"101111000001110001110100001011001000",--18894
"111110001110001001000011100000000000",--18895
"101111000001110010000100000110101000",--18896
"111110010000000001100011000000000000",--18897
"111110001100011000000011000000000000",--18898
"111110001110001001100011000000000000",--18899
"101111000001110001110100001010100010",--18900
"111110001110001001000011100000000000",--18901
"101111000001110010000100000110011000",--18902
"111110010000000001100011000000000000",--18903
"111110001100011000000011000000000000",--18904
"111110001110001001100011000000000000",--18905
"101111000001110001110100001010000000",--18906
"111110001110001001000011100000000000",--18907
"101111000001110010000100000110001000",--18908
"111110010000000001100011000000000000",--18909
"111110001100011000000011000000000000",--18910
"111110001110001001100011000000000000",--18911
"101111000001110001110100001001000100",--18912
"111110001110001001000011100000000000",--18913
"101111000001110010000100000101110000",--18914
"111110010000000001100011000000000000",--18915
"111110001100011000000011000000000000",--18916
"111110001110001001100011000000000000",--18917
"101111000001110001110100001000010000",--18918
"111110001110001001000011100000000000",--18919
"101111000001110010000100000101010000",--18920
"111110010000000001100011000000000000",--18921
"111110001100011000000011000000000000",--18922
"111110001110001001100011000000000000",--18923
"101111000001110001110100000111001000",--18924
"111110001110001001000011100000000000",--18925
"101111000001110010000100000100110000",--18926
"111110010000000001100011000000000000",--18927
"111110001100011000000011000000000000",--18928
"111110001110001001100011000000000000",--18929
"101111000001110001110100000110000000",--18930
"111110001110001001000011100000000000",--18931
"101111000001110010000100000100010000",--18932
"111110010000000001100011000000000000",--18933
"111110001100011000000011000000000000",--18934
"111110001110001001100011000000000000",--18935
"101111000001110001110100000100010000",--18936
"111110001110001001000011100000000000",--18937
"101111000001110010000100000011100000",--18938
"111110010000000001100011000000000000",--18939
"111110001100011000000011000000000000",--18940
"111110001110001001100011000000000000",--18941
"101111000001110010000100000010000000",--18942
"111110010000001001000100000000000000",--18943
"101111000001110010010100000010100000",--18944
"111110010010000001100011000000000000",--18945
"111110001100011000000011000000000000",--18946
"111110010000001001100011000000000000",--18947
"001001111100000001001111111111110100",--18948
"001011111100000000111111111111110011",--18949
"101110001101111000000010100000000000",--18950
"101110000011111000000001100000000000",--18951
"001001111100000111111111111111110010",--18952
"101001111100010111100000000000001111",--18953
"000111000000000000000000001101001100",--18954
"101001111100000111100000000000001111",--18955
"001101111100000111111111111111110010",--18956
"111110000110000000010001100000000000",--18957
"111110000110011000000001100000000000",--18958
"001111111100000001001111111111110011",--18959
"111110001000001000110001100000000000",--18960
"001101111100000000011111111111110100",--18961
"010100000011000000000000000000000100",--18962
"101111001001110001000011111111001001",--18963
"101111001001100001000000111111011010",--18964
"111110001000010000110001100000000000",--18965
"000101000000000000000100101000011011",--18966
"011000000011000000000000000000000011",--18967
"101111001001110001001011111111001001",--18968
"101111001001100001000000111111011010",--18969
"111110001000010000110001100000000000",--18970
"101111000001110001000100000111110000",--18971
"111110000110001001000001100000000000",--18972
"101111001001110001000011111010100010",--18973
"101111001001100001001111100110000010",--18974
"111110000110001001000001100000000000",--18975
"101110000110110000000010000000000000",--18976
"111110000110010001000001100000000000",--18977
"001111111100000001001111111111110101",--18978
"101110001001111000000010100000000001",--18979
"101111001101110001100011100011010001",--18980
"101111001101100001101011011100010111",--18981
"001011111100000000111111111111110100",--18982
"010110001101000001010000000000000010",--18983
"101111000001110000110100000101110000",--18984
"000101000000000000000100101010010110",--18985
"001111000000000001010000000100101011",--18986
"001101111100000000011111111111110110",--18987
"001111000010000001100000000000000001",--18988
"111110001010010001100010100000000000",--18989
"001101111100000000011111111111110111",--18990
"001111000010000001100000000000000001",--18991
"111110001100100000000011000000000000",--18992
"111110001010001001100010100000000000",--18993
"111110001000011000000010000000000000",--18994
"111110001010001001000010000000000001",--18995
"010110001001000000010000000000000010",--18996
"101001000000000000010000000000000001",--18997
"000101000000000000000100101000111100",--18998
"011010001001000000100000000000000010",--18999
"101001000000000000011111111111111111",--19000
"000101000000000000000100101000111100",--19001
"101000000001111000000000100000000000",--19002
"000101000000000000000100101000111101",--19003
"111110001000011000000010000000000000",--19004
"111110001000001001000010100000000000",--19005
"101111000001110001100100001011110010",--19006
"111110001100001001010011000000000000",--19007
"101111001111110001110011110100110010",--19008
"101111001111100001110001011001000011",--19009
"111110001100001001110011000000000000",--19010
"101111000001110001110100001011001000",--19011
"111110001110001001010011100000000000",--19012
"101111000001110010000100000110101000",--19013
"111110010000000001100011000000000000",--19014
"111110001100011000000011000000000000",--19015
"111110001110001001100011000000000000",--19016
"101111000001110001110100001010100010",--19017
"111110001110001001010011100000000000",--19018
"101111000001110010000100000110011000",--19019
"111110010000000001100011000000000000",--19020
"111110001100011000000011000000000000",--19021
"111110001110001001100011000000000000",--19022
"101111000001110001110100001010000000",--19023
"111110001110001001010011100000000000",--19024
"101111000001110010000100000110001000",--19025
"111110010000000001100011000000000000",--19026
"111110001100011000000011000000000000",--19027
"111110001110001001100011000000000000",--19028
"101111000001110001110100001001000100",--19029
"111110001110001001010011100000000000",--19030
"101111000001110010000100000101110000",--19031
"111110010000000001100011000000000000",--19032
"111110001100011000000011000000000000",--19033
"111110001110001001100011000000000000",--19034
"101111000001110001110100001000010000",--19035
"111110001110001001010011100000000000",--19036
"101111000001110010000100000101010000",--19037
"111110010000000001100011000000000000",--19038
"111110001100011000000011000000000000",--19039
"111110001110001001100011000000000000",--19040
"101111000001110001110100000111001000",--19041
"111110001110001001010011100000000000",--19042
"101111000001110010000100000100110000",--19043
"111110010000000001100011000000000000",--19044
"111110001100011000000011000000000000",--19045
"111110001110001001100011000000000000",--19046
"101111000001110001110100000110000000",--19047
"111110001110001001010011100000000000",--19048
"101111000001110010000100000100010000",--19049
"111110010000000001100011000000000000",--19050
"111110001100011000000011000000000000",--19051
"111110001110001001100011000000000000",--19052
"101111000001110001110100000100010000",--19053
"111110001110001001010011100000000000",--19054
"101111000001110010000100000011100000",--19055
"111110010000000001100011000000000000",--19056
"111110001100011000000011000000000000",--19057
"111110001110001001100011000000000000",--19058
"101111000001110010000100000010000000",--19059
"111110010000001001010100000000000000",--19060
"101111000001110010010100000010100000",--19061
"111110010010000001100011000000000000",--19062
"111110001100011000000011000000000000",--19063
"111110010000001001100011000000000000",--19064
"001001111100000000011111111111110011",--19065
"001011111100000001001111111111110010",--19066
"101110001011111000000010000000000000",--19067
"101110000011111000000001100000000000",--19068
"101110001101111000000010100000000000",--19069
"001001111100000111111111111111110001",--19070
"101001111100010111100000000000010000",--19071
"000111000000000000000000001101001100",--19072
"101001111100000111100000000000010000",--19073
"001101111100000111111111111111110001",--19074
"111110000110000000010001100000000000",--19075
"111110000110011000000001100000000000",--19076
"001111111100000001001111111111110010",--19077
"111110001000001000110001100000000000",--19078
"001101111100000000011111111111110011",--19079
"010100000011000000000000000000000100",--19080
"101111001001110001000011111111001001",--19081
"101111001001100001000000111111011010",--19082
"111110001000010000110001100000000000",--19083
"000101000000000000000100101010010001",--19084
"011000000011000000000000000000000011",--19085
"101111001001110001001011111111001001",--19086
"101111001001100001000000111111011010",--19087
"111110001000010000110001100000000000",--19088
"101111000001110001000100000111110000",--19089
"111110000110001001000001100000000000",--19090
"101111001001110001000011111010100010",--19091
"101111001001100001001111100110000010",--19092
"111110000110001001000001100000000000",--19093
"101110000110110000000010000000000000",--19094
"111110000110010001000001100000000000",--19095
"101111001001110001000011111000011001",--19096
"101111001001100001001001100110011010",--19097
"101111000001110001010011111100000000",--19098
"001111111100000001101111111111110100",--19099
"111110001010010001100010100000000000",--19100
"111110001010001001010010100000000000",--19101
"111110001000010001010010000000000000",--19102
"101111000001110001010011111100000000",--19103
"111110001010010000110001100000000000",--19104
"111110000110001000110001100000000000",--19105
"111110001000010000110001100000000000",--19106
"011010000111000000000000000000000001",--19107
"101110000001111000000001100000000000",--19108
"101111000001110001000100001101111111",--19109
"111110001000001000110001100000000000",--19110
"101111001001110001000100000001010101",--19111
"101111001001100001000101010101010101",--19112
"111110000110001001000001100000000000",--19113
"001011000000000000110000000100100101",--19114
"001101000000000000100000000100110000",--19115
"001101000100000000010000000000000000",--19116
"001101000010000000110000000000000000",--19117
"010011000111000000000000000010110100",--19118
"001001111100000000011111111111110111",--19119
"001001111100000000101111111111110110",--19120
"010011000111011000110000000010100010",--19121
"001101000110000001000000000101101101",--19122
"001111000000000000110000000100101010",--19123
"001101001000000001010000000000000101",--19124
"001111001010000001000000000000000000",--19125
"111110000110010001000001100000000000",--19126
"001111000000000001000000000100101011",--19127
"001111001010000001010000000000000001",--19128
"111110001000010001010010000000000000",--19129
"001111000000000001010000000100101100",--19130
"001111001010000001100000000000000010",--19131
"111110001010010001100010100000000000",--19132
"001101000110000000110000000010111110",--19133
"001101001000000001010000000000000001",--19134
"011111001011000000010000000000110111",--19135
"001111000110000001100000000000000000",--19136
"111110001100010000110011000000000000",--19137
"001111000110000001110000000000000001",--19138
"111110001100001001110011000000000000",--19139
"001111000000000001110000000011111011",--19140
"111110001100001001110011100000000000",--19141
"111110001110000001000011100000000001",--19142
"001101001000000001000000000000000100",--19143
"001111001000000010000000000000000001",--19144
"010110010001000001110000000000000111",--19145
"001111000000000001110000000011111100",--19146
"111110001100001001110011100000000000",--19147
"111110001110000001010011100000000001",--19148
"001111001000000010000000000000000010",--19149
"010110010001000001110000000000000010",--19150
"001111000110000001110000000000000001",--19151
"011110001111000000000000000000100100",--19152
"001111000110000001100000000000000010",--19153
"111110001100010001000011000000000000",--19154
"001111000110000001110000000000000011",--19155
"111110001100001001110011000000000000",--19156
"001111000000000001110000000011111010",--19157
"111110001100001001110011100000000000",--19158
"111110001110000000110011100000000001",--19159
"001111001000000010000000000000000000",--19160
"010110010001000001110000000000000111",--19161
"001111000000000001110000000011111100",--19162
"111110001100001001110011100000000000",--19163
"111110001110000001010011100000000001",--19164
"001111001000000010000000000000000010",--19165
"010110010001000001110000000000000010",--19166
"001111000110000001110000000000000011",--19167
"011110001111000000000000000000010010",--19168
"001111000110000001100000000000000100",--19169
"111110001100010001010010100000000000",--19170
"001111000110000001100000000000000101",--19171
"111110001010001001100010100000000000",--19172
"001111000000000001100000000011111010",--19173
"111110001010001001100011000000000000",--19174
"111110001100000000110001100000000001",--19175
"001111001000000001100000000000000000",--19176
"010110001101000000110000000001100001",--19177
"001111000000000000110000000011111011",--19178
"111110001010001000110001100000000000",--19179
"111110000110000001000001100000000001",--19180
"001111001000000001000000000000000001",--19181
"010110001001000000110000000001011100",--19182
"001111000110000000110000000000000101",--19183
"010010000111000000000000000001011010",--19184
"001011000000000001010000000100101111",--19185
"000101000000000000000100101100111111",--19186
"001011000000000001100000000100101111",--19187
"000101000000000000000100101100111111",--19188
"001011000000000001100000000100101111",--19189
"000101000000000000000100101100111111",--19190
"011111001011000000100000000000001100",--19191
"001111000110000001100000000000000000",--19192
"011010001101000000000000000001010001",--19193
"001111000110000001100000000000000001",--19194
"111110001100001000110001100000000000",--19195
"001111000110000001100000000000000010",--19196
"111110001100001001000010000000000000",--19197
"111110000110000001000001100000000000",--19198
"001111000110000001000000000000000011",--19199
"111110001000001001010010000000000000",--19200
"111110000110000001000001100000000000",--19201
"001011000000000000110000000100101111",--19202
"000101000000000000000100101100111111",--19203
"001111000110000001100000000000000000",--19204
"010010001101000000000000000001000101",--19205
"001111000110000001110000000000000001",--19206
"111110001110001000110011100000000000",--19207
"001111000110000010000000000000000010",--19208
"111110010000001001000100000000000000",--19209
"111110001110000010000011100000000000",--19210
"001111000110000010000000000000000011",--19211
"111110010000001001010100000000000000",--19212
"111110001110000010000011100000000000",--19213
"111110000110001000110100000000000000",--19214
"001101001000000001100000000000000100",--19215
"001111001100000010010000000000000000",--19216
"111110010000001010010100000000000000",--19217
"111110001000001001000100100000000000",--19218
"001111001100000010100000000000000001",--19219
"111110010010001010100100100000000000",--19220
"111110010000000010010100000000000000",--19221
"111110001010001001010100100000000000",--19222
"001111001100000010100000000000000010",--19223
"111110010010001010100100100000000000",--19224
"111110010000000010010100000000000000",--19225
"001101001000000001100000000000000011",--19226
"011100001101000000000000000000000011",--19227
"101110010001111000000001100000000000",--19228
"011111001011000000110000000000010000",--19229
"000101000000000000000100101100101101",--19230
"111110001000001001010100100000000000",--19231
"001101001000000001100000000000001001",--19232
"001111001100000010100000000000000000",--19233
"111110010010001010100100100000000000",--19234
"111110010000000010010100000000000000",--19235
"111110001010001000110010100000000000",--19236
"001111001100000010010000000000000001",--19237
"111110001010001010010010100000000000",--19238
"111110010000000001010010100000000000",--19239
"111110000110001001000001100000000000",--19240
"001111001100000001000000000000000010",--19241
"111110000110001001000001100000000000",--19242
"111110001010000000110001100000000000",--19243
"011111001011000000110000000000000001",--19244
"111110000110010000010001100000000000",--19245
"111110001110001001110010000000000000",--19246
"111110001100001000110001100000000000",--19247
"111110001000010000110001100000000000",--19248
"010110000111000000000000000000011001",--19249
"001101001000000001000000000000000110",--19250
"011100001001000000000000000000000110",--19251
"111110000110100000000001100000000000",--19252
"111110001110010000110001100000000000",--19253
"001111000110000001000000000000000100",--19254
"111110000110001001000001100000000000",--19255
"001011000000000000110000000100101111",--19256
"000101000000000000000100101100111111",--19257
"111110000110100000000001100000000000",--19258
"111110001110000000110001100000000000",--19259
"001111000110000001000000000000000100",--19260
"111110000110001001000001100000000000",--19261
"001011000000000000110000000100101111",--19262
"001111000000000000110000000100101111",--19263
"101111001001110001001011110111001100",--19264
"101111001001100001001100110011001101",--19265
"010110001001000000110000000000001000",--19266
"101000000011111000000001000000000000",--19267
"101001000000000000010000000000000001",--19268
"001001111100000111111111111111110101",--19269
"101001111100010111100000000000001100",--19270
"000111000000000000000000110101111110",--19271
"101001111100000111100000000000001100",--19272
"001101111100000111111111111111110101",--19273
"011100000011000000000000000000001001",--19274
"101001000000000000010000000000000001",--19275
"001101111100000000101111111111110110",--19276
"001001111100000111111111111111110101",--19277
"101001111100010111100000000000001100",--19278
"000111000000000000000000111111111011",--19279
"101001111100000111100000000000001100",--19280
"001101111100000111111111111111110101",--19281
"011100000011000000000000000000110110",--19282
"000101000000000000000100101101100011",--19283
"101001000000000000010000000000000001",--19284
"001101111100000000101111111111110111",--19285
"001001111100000111111111111111110101",--19286
"101001111100010111100000000000001100",--19287
"000111000000000000000000110101111110",--19288
"101001111100000111100000000000001100",--19289
"001101111100000111111111111111110101",--19290
"011100000011000000000000000000101101",--19291
"101001000000000000010000000000000001",--19292
"001101111100000000101111111111110110",--19293
"101001111100010111100000000000001100",--19294
"000111000000000000000000111111111011",--19295
"101001111100000111100000000000001100",--19296
"001101111100000111111111111111110101",--19297
"011100000011000000000000000000100110",--19298
"101111000111110000110011101111011010",--19299
"101111000111100000110111010000001101",--19300
"001111111100000001001111111111111010",--19301
"111110001000001000110001100000000000",--19302
"001111000000000001000000000100100110",--19303
"001111000000000001010000000101100100",--19304
"111110001000001001010010000000000000",--19305
"001111000000000001010000000100100111",--19306
"001111000000000001100000000101100101",--19307
"111110001010001001100010100000000000",--19308
"111110001000000001010010000000000000",--19309
"001111000000000001010000000100101000",--19310
"001111000000000001100000000101100110",--19311
"111110001010001001100010100000000000",--19312
"111110001000000001010010000000000010",--19313
"010110001001000000000000000000000001",--19314
"000101000000000000000100101101110101",--19315
"101110000001111000000010000000000000",--19316
"111110000110001001000001100000000000",--19317
"001101111100000000011111111111111000",--19318
"001101000010000000010000000000000111",--19319
"001111000010000001000000000000000000",--19320
"111110000110001001000001100000000000",--19321
"001111000000000001000000000100100000",--19322
"001111000000000001010000000100100011",--19323
"111110000110001001010010100000000000",--19324
"111110001000000001010010000000000000",--19325
"001011000000000001000000000100100000",--19326
"001111000000000001000000000100100001",--19327
"001111000000000001010000000100100100",--19328
"111110000110001001010010100000000000",--19329
"111110001000000001010010000000000000",--19330
"001011000000000001000000000100100001",--19331
"001111000000000001000000000100100010",--19332
"001111000000000001010000000100100101",--19333
"111110000110001001010001100000000000",--19334
"111110001000000000110001100000000000",--19335
"001011000000000000110000000100100010",--19336
"001101111100000000011111111111111011",--19337
"101001000010010001000000000000000010",--19338
"001101111100000000011111111111111110",--19339
"001101111100000000101111111111111111",--19340
"001101111100000000110000000000000000",--19341
"010111001000000000001111100000000000",--19342
"000101000000000000000100000011011011",--19343
"001111000110000000110000000000000000",--19344
"001011000000000000110000000100010010",--19345
"001111000110000000110000000000000001",--19346
"001011000000000000110000000100010011",--19347
"001111000110000000110000000000000010",--19348
"001011000000000000110000000100010100",--19349
"001101000000000001000000000110101010",--19350
"101001001000010001000000000000000001",--19351
"001001111100000000110000000000000000",--19352
"001001111100000000101111111111111111",--19353
"001001111100000000011111111111111110",--19354
"010111001001000000000000000010010001",--19355
"001101001000000001010000000101101101",--19356
"001101001010000001100000000000001010",--19357
"001101001010000001110000000000000001",--19358
"001111000110000000110000000000000000",--19359
"001101001010000010000000000000000101",--19360
"001111010000000001000000000000000000",--19361
"111110000110010001000001100000000000",--19362
"001011001100000000110000000000000000",--19363
"001111000110000000110000000000000001",--19364
"001111010000000001000000000000000001",--19365
"111110000110010001000001100000000000",--19366
"001011001100000000110000000000000001",--19367
"001111000110000000110000000000000010",--19368
"001111010000000001000000000000000010",--19369
"111110000110010001000001100000000000",--19370
"001011001100000000110000000000000010",--19371
"011111001111000000100000000000001110",--19372
"001101001010000001010000000000000100",--19373
"001111001100000000110000000000000000",--19374
"001111001100000001000000000000000001",--19375
"001111001100000001010000000000000010",--19376
"001111001010000001100000000000000000",--19377
"111110001100001000110001100000000000",--19378
"001111001010000001100000000000000001",--19379
"111110001100001001000010000000000000",--19380
"111110000110000001000001100000000000",--19381
"001111001010000001000000000000000010",--19382
"111110001000001001010010000000000000",--19383
"111110000110000001000001100000000000",--19384
"001011001100000000110000000000000011",--19385
"000101000000000000000100101111100000",--19386
"010111001111000000100000000000100100",--19387
"001111001100000000110000000000000000",--19388
"001111001100000001000000000000000001",--19389
"001111001100000001010000000000000010",--19390
"111110000110001000110011000000000000",--19391
"001101001010000010000000000000000100",--19392
"001111010000000001110000000000000000",--19393
"111110001100001001110011000000000000",--19394
"111110001000001001000011100000000000",--19395
"001111010000000010000000000000000001",--19396
"111110001110001010000011100000000000",--19397
"111110001100000001110011000000000000",--19398
"111110001010001001010011100000000000",--19399
"001111010000000010000000000000000010",--19400
"111110001110001010000011100000000000",--19401
"111110001100000001110011000000000000",--19402
"001101001010000010000000000000000011",--19403
"011100010001000000000000000000000011",--19404
"101110001101111000000001100000000000",--19405
"011111001111000000110000000000010000",--19406
"000101000000000000000100101111011110",--19407
"111110001000001001010011100000000000",--19408
"001101001010000001010000000000001001",--19409
"001111001010000010000000000000000000",--19410
"111110001110001010000011100000000000",--19411
"111110001100000001110011000000000000",--19412
"111110001010001000110010100000000000",--19413
"001111001010000001110000000000000001",--19414
"111110001010001001110010100000000000",--19415
"111110001100000001010010100000000000",--19416
"111110000110001001000001100000000000",--19417
"001111001010000001000000000000000010",--19418
"111110000110001001000001100000000000",--19419
"111110001010000000110001100000000000",--19420
"011111001111000000110000000000000001",--19421
"111110000110010000010001100000000000",--19422
"001011001100000000110000000000000011",--19423
"101001001000010001000000000000000001",--19424
"010111001001000000000000000001001011",--19425
"001101001000000001010000000101101101",--19426
"001101001010000001100000000000001010",--19427
"001101001010000001110000000000000001",--19428
"001111000110000000110000000000000000",--19429
"001101001010000010000000000000000101",--19430
"001111010000000001000000000000000000",--19431
"111110000110010001000001100000000000",--19432
"001011001100000000110000000000000000",--19433
"001111000110000000110000000000000001",--19434
"001111010000000001000000000000000001",--19435
"111110000110010001000001100000000000",--19436
"001011001100000000110000000000000001",--19437
"001111000110000000110000000000000010",--19438
"001111010000000001000000000000000010",--19439
"111110000110010001000001100000000000",--19440
"001011001100000000110000000000000010",--19441
"011111001111000000100000000000001110",--19442
"001101001010000001010000000000000100",--19443
"001111001100000000110000000000000000",--19444
"001111001100000001000000000000000001",--19445
"001111001100000001010000000000000010",--19446
"001111001010000001100000000000000000",--19447
"111110001100001000110001100000000000",--19448
"001111001010000001100000000000000001",--19449
"111110001100001001000010000000000000",--19450
"111110000110000001000001100000000000",--19451
"001111001010000001000000000000000010",--19452
"111110001000001001010010000000000000",--19453
"111110000110000001000001100000000000",--19454
"001011001100000000110000000000000011",--19455
"000101000000000000000100110000100110",--19456
"010111001111000000100000000000100100",--19457
"001111001100000000110000000000000000",--19458
"001111001100000001000000000000000001",--19459
"001111001100000001010000000000000010",--19460
"111110000110001000110011000000000000",--19461
"001101001010000010000000000000000100",--19462
"001111010000000001110000000000000000",--19463
"111110001100001001110011000000000000",--19464
"111110001000001001000011100000000000",--19465
"001111010000000010000000000000000001",--19466
"111110001110001010000011100000000000",--19467
"111110001100000001110011000000000000",--19468
"111110001010001001010011100000000000",--19469
"001111010000000010000000000000000010",--19470
"111110001110001010000011100000000000",--19471
"111110001100000001110011000000000000",--19472
"001101001010000010000000000000000011",--19473
"011100010001000000000000000000000011",--19474
"101110001101111000000001100000000000",--19475
"011111001111000000110000000000010000",--19476
"000101000000000000000100110000100100",--19477
"111110001000001001010011100000000000",--19478
"001101001010000001010000000000001001",--19479
"001111001010000010000000000000000000",--19480
"111110001110001010000011100000000000",--19481
"111110001100000001110011000000000000",--19482
"111110001010001000110010100000000000",--19483
"001111001010000001110000000000000001",--19484
"111110001010001001110010100000000000",--19485
"111110001100000001010010100000000000",--19486
"111110000110001001000001100000000000",--19487
"001111001010000001000000000000000010",--19488
"111110000110001001000001100000000000",--19489
"111110001010000000110001100000000000",--19490
"011111001111000000110000000000000001",--19491
"111110000110010000010001100000000000",--19492
"001011001100000000110000000000000011",--19493
"101001001000010000100000000000000001",--19494
"101000000111111000000000100000000000",--19495
"001001111100000111111111111111111101",--19496
"101001111100010111100000000000000100",--19497
"000111000000000000000000011001101110",--19498
"101001111100000111100000000000000100",--19499
"001101111100000111111111111111111101",--19500
"001101111100000000011111111111111110",--19501
"001101000010000000100000000001110110",--19502
"001101000100000000100000000000000000",--19503
"001111000100000000110000000000000000",--19504
"001101111100000000111111111111111111",--19505
"001111000110000001000000000000000000",--19506
"111110000110001001000001100000000000",--19507
"001111000100000001000000000000000001",--19508
"001111000110000001010000000000000001",--19509
"111110001000001001010010000000000000",--19510
"111110000110000001000001100000000000",--19511
"001111000100000001000000000000000010",--19512
"001111000110000001010000000000000010",--19513
"111110001000001001010010000000000000",--19514
"111110000110000001000001100000000000",--19515
"011010000111000000000000001011000110",--19516
"001101000010000000110000000001110111",--19517
"101111001001110001000100111001101110",--19518
"101111001001100001000110101100101000",--19519
"001011000000000001000000000100101101",--19520
"001101000000000000100000000100110000",--19521
"001011111100000000111111111111111101",--19522
"001001111100000000111111111111111100",--19523
"101000000001111000000000100000000000",--19524
"001001111100000111111111111111111011",--19525
"101001111100010111100000000000000110",--19526
"000111000000000000000010110111111111",--19527
"101001111100000111100000000000000110",--19528
"001101111100000111111111111111111011",--19529
"001111000000000000110000000100101101",--19530
"101111001001110001001011110111001100",--19531
"101111001001100001001100110011001101",--19532
"010110000111000001000000010101111010",--19533
"101111001001110001000100110010111110",--19534
"101111001001100001001011110000100000",--19535
"010110001001000000110000010101110111",--19536
"001101000000000000010000000100101001",--19537
"001101000010000000010000000101101101",--19538
"001101000010000000100000000000000001",--19539
"011111000101000000010000000000010011",--19540
"001101111100000000101111111111111100",--19541
"001101000100000000100000000000000000",--19542
"001101000000000000110000000100101110",--19543
"001011000000000000000000000100100110",--19544
"001011000000000000000000000100100111",--19545
"001011000000000000000000000100101000",--19546
"101001000110010001000000000000000001",--19547
"101001000110010000110000000000000001",--19548
"001110000100000000110001100000000000",--19549
"011110000111000000000000000000000010",--19550
"101110000001111000000001100000000000",--19551
"000101000000000000000100110001100101",--19552
"010110000111000000000000000000000010",--19553
"101110000011111000000001100000000000",--19554
"000101000000000000000100110001100101",--19555
"101110000101111000000001100000000000",--19556
"101110000111111000000001100000000010",--19557
"001011001000000000110000000100100110",--19558
"000101000000000000000100110010111110",--19559
"011111000101000000100000000000001000",--19560
"001101000010000000100000000000000100",--19561
"001111000100010000110000000000000000",--19562
"001011000000000000110000000100100110",--19563
"001111000100010000110000000000000001",--19564
"001011000000000000110000000100100111",--19565
"001111000100010000110000000000000010",--19566
"001011000000000000110000000100101000",--19567
"000101000000000000000100110010111110",--19568
"001111000000000000110000000100101010",--19569
"001101000010000000100000000000000101",--19570
"001111000100000001000000000000000000",--19571
"111110000110010001000001100000000000",--19572
"001111000000000001000000000100101011",--19573
"001111000100000001010000000000000001",--19574
"111110001000010001010010000000000000",--19575
"001111000000000001010000000100101100",--19576
"001111000100000001100000000000000010",--19577
"111110001010010001100010100000000000",--19578
"001101000010000000100000000000000100",--19579
"001111000100000001100000000000000000",--19580
"111110000110001001100011000000000000",--19581
"001111000100000001110000000000000001",--19582
"111110001000001001110011100000000000",--19583
"001111000100000010000000000000000010",--19584
"111110001010001010000100000000000000",--19585
"001101000010000000100000000000000011",--19586
"011100000101000000000000000000000100",--19587
"001011000000000001100000000100100110",--19588
"001011000000000001110000000100100111",--19589
"001011000000000010000000000100101000",--19590
"000101000000000000000100110010100100",--19591
"001101000010000000100000000000001001",--19592
"001111000100000010010000000000000010",--19593
"111110001000001010010100100000000000",--19594
"001111000100000010100000000000000001",--19595
"111110001010001010100101000000000000",--19596
"111110010010000010100100100000000000",--19597
"101111000001110010100011111100000000",--19598
"111110010010001010100100100000000000",--19599
"111110001100000010010011000000000000",--19600
"001011000000000001100000000100100110",--19601
"001111000100000001100000000000000010",--19602
"111110000110001001100011000000000000",--19603
"001111000100000010010000000000000000",--19604
"111110001010001010010010100000000000",--19605
"111110001100000001010010100000000000",--19606
"101111000001110001100011111100000000",--19607
"111110001010001001100010100000000000",--19608
"111110001110000001010010100000000000",--19609
"001011000000000001010000000100100111",--19610
"001111000100000001010000000000000001",--19611
"111110000110001001010001100000000000",--19612
"001111000100000001010000000000000000",--19613
"111110001000001001010010000000000000",--19614
"111110000110000001000001100000000000",--19615
"101111000001110001000011111100000000",--19616
"111110000110001001000001100000000000",--19617
"111110010000000000110001100000000000",--19618
"001011000000000000110000000100101000",--19619
"001111000000000000110000000100100110",--19620
"111110000110001000110001100000000000",--19621
"001111000000000001000000000100100111",--19622
"111110001000001001000010000000000000",--19623
"111110000110000001000001100000000000",--19624
"001111000000000001000000000100101000",--19625
"111110001000001001000010000000000000",--19626
"111110000110000001000001100000000000",--19627
"111110000110100000000001100000000000",--19628
"011110000111000000000000000000000010",--19629
"101110000011111000000001100000000000",--19630
"000101000000000000000100110010110101",--19631
"001101000010000000100000000000000110",--19632
"011100000101000000000000000000000010",--19633
"111110000110011000000001100000000000",--19634
"000101000000000000000100110010110101",--19635
"111110000110011000000001100000000010",--19636
"001111000000000001000000000100100110",--19637
"111110001000001000110010000000000000",--19638
"001011000000000001000000000100100110",--19639
"001111000000000001000000000100100111",--19640
"111110001000001000110010000000000000",--19641
"001011000000000001000000000100100111",--19642
"001111000000000001000000000100101000",--19643
"111110001000001000110001100000000000",--19644
"001011000000000000110000000100101000",--19645
"001101000010000000100000000000000000",--19646
"001101000010000000110000000000001000",--19647
"001111000110000000110000000000000000",--19648
"001011000000000000110000000100100011",--19649
"001111000110000000110000000000000001",--19650
"001011000000000000110000000100100100",--19651
"001111000110000000110000000000000010",--19652
"001011000000000000110000000100100101",--19653
"001001111100000000011111111111111011",--19654
"011111000101000000010000000000100011",--19655
"001111000000000000110000000100101010",--19656
"001101000010000000100000000000000101",--19657
"001111000100000001000000000000000000",--19658
"111110000110010001000001100000000000",--19659
"101111001001110001000011110101001100",--19660
"101111001001100001001100110011001101",--19661
"111110000110001001000010000000000000",--19662
"101110001000110000000010000000000000",--19663
"101111000001110001010100000110100000",--19664
"111110001000001001010010000000000000",--19665
"111110000110010001000001100000000000",--19666
"101111000001110001000100000100100000",--19667
"001111000000000001010000000100101100",--19668
"001111000100000001100000000000000010",--19669
"111110001010010001100010100000000000",--19670
"101111001101110001100011110101001100",--19671
"101111001101100001101100110011001101",--19672
"111110001010001001100011000000000000",--19673
"101110001100110000000011000000000000",--19674
"101111000001110001110100000110100000",--19675
"111110001100001001110011000000000000",--19676
"111110001010010001100010100000000000",--19677
"101111000001110001100100000100100000",--19678
"010110001001000000110000000000000101",--19679
"010110001101000001010000000000000010",--19680
"101111000001110000110100001101111111",--19681
"000101000000000000000100110011101001",--19682
"101110000001111000000001100000000000",--19683
"000101000000000000000100110011101001",--19684
"010110001101000001010000000000000010",--19685
"101110000001111000000001100000000000",--19686
"000101000000000000000100110011101001",--19687
"101111000001110000110100001101111111",--19688
"001011000000000000110000000100100100",--19689
"000101000000000000000100111000100100",--19690
"011111000101000000100000000000001111",--19691
"001111000000000000110000000100101011",--19692
"101111000001110001000011111010000000",--19693
"111110000110001001000001100000000000",--19694
"001001111100000111111111111111111010",--19695
"000111000000000000000111011000000010",--19696
"001101111100000111111111111111111010",--19697
"111110000110001000110001100000000000",--19698
"101111000001110001000100001101111111",--19699
"111110001000001000110010000000000000",--19700
"001011000000000001000000000100100011",--19701
"101111000001110001000100001101111111",--19702
"111110000110010000010001100000000010",--19703
"111110001000001000110001100000000000",--19704
"001011000000000000110000000100100100",--19705
"000101000000000000000100111000100100",--19706
"011111000101000000110000000000011111",--19707
"001111000000000000110000000100101010",--19708
"001101000010000000100000000000000101",--19709
"001111000100000001000000000000000000",--19710
"111110000110010001000001100000000000",--19711
"001111000000000001000000000100101100",--19712
"001111000100000001010000000000000010",--19713
"111110001000010001010010000000000000",--19714
"111110000110001000110001100000000000",--19715
"111110001000001001000010000000000000",--19716
"111110000110000001000001100000000000",--19717
"111110000110100000000001100000000000",--19718
"101111001001110001000011110111001100",--19719
"101111001001100001001100110011001100",--19720
"111110000110001001000001100000000000",--19721
"101110000110110000000010000000000000",--19722
"111110000110010001000001100000000000",--19723
"101111001001110001000100000001001001",--19724
"101111001001100001000000111111011011",--19725
"111110000110001001000001100000000000",--19726
"001001111100000111111111111111111010",--19727
"000111000000000000000111010110111000",--19728
"001101111100000111111111111111111010",--19729
"111110000110001000110001100000000000",--19730
"101111000001110001000100001101111111",--19731
"111110000110001001000010000000000000",--19732
"001011000000000001000000000100100100",--19733
"111110000110010000010001100000000010",--19734
"101111000001110001000100001101111111",--19735
"111110000110001001000001100000000000",--19736
"001011000000000000110000000100100101",--19737
"000101000000000000000100111000100100",--19738
"011111000101000001000000000100001000",--19739
"001111000000000000110000000100101010",--19740
"001101000010000000100000000000000101",--19741
"001111000100000001000000000000000000",--19742
"111110000110010001000001100000000000",--19743
"001101000010000000110000000000000100",--19744
"001111000110000001000000000000000000",--19745
"111110001000100000000010000000000000",--19746
"111110000110001001000001100000000000",--19747
"001111000000000001000000000100101100",--19748
"001111000100000001010000000000000010",--19749
"111110001000010001010010000000000000",--19750
"001111000110000001010000000000000010",--19751
"111110001010100000000010100000000000",--19752
"111110001000001001010010000000000000",--19753
"111110000110001000110010100000000000",--19754
"111110001000001001000011000000000000",--19755
"111110001010000001100010100000000000",--19756
"101110000111111000000011000000000001",--19757
"101111001111110001110011100011010001",--19758
"101111001111100001111011011100010111",--19759
"001001111100000000111111111111111010",--19760
"001001111100000000101111111111111001",--19761
"001011111100000001011111111111111000",--19762
"010110001111000001100000000000000010",--19763
"101111000001110000110100000101110000",--19764
"000101000000000000000100110110011001",--19765
"111110000110011000000001100000000000",--19766
"111110001000001000110001100000000001",--19767
"010110000111000000010000000000000010",--19768
"101001000000000001000000000000000001",--19769
"000101000000000000000100110101000000",--19770
"011010000111000000100000000000000010",--19771
"101001000000000001001111111111111111",--19772
"000101000000000000000100110101000000",--19773
"101000000001111000000010000000000000",--19774
"000101000000000000000100110101000001",--19775
"111110000110011000000001100000000000",--19776
"111110000110001000110010000000000000",--19777
"101111000001110001100100001011110010",--19778
"111110001100001001000011000000000000",--19779
"101111001111110001110011110100110010",--19780
"101111001111100001110001011001000011",--19781
"111110001100001001110011000000000000",--19782
"101111000001110001110100001011001000",--19783
"111110001110001001000011100000000000",--19784
"101111000001110010000100000110101000",--19785
"111110010000000001100011000000000000",--19786
"111110001100011000000011000000000000",--19787
"111110001110001001100011000000000000",--19788
"101111000001110001110100001010100010",--19789
"111110001110001001000011100000000000",--19790
"101111000001110010000100000110011000",--19791
"111110010000000001100011000000000000",--19792
"111110001100011000000011000000000000",--19793
"111110001110001001100011000000000000",--19794
"101111000001110001110100001010000000",--19795
"111110001110001001000011100000000000",--19796
"101111000001110010000100000110001000",--19797
"111110010000000001100011000000000000",--19798
"111110001100011000000011000000000000",--19799
"111110001110001001100011000000000000",--19800
"101111000001110001110100001001000100",--19801
"111110001110001001000011100000000000",--19802
"101111000001110010000100000101110000",--19803
"111110010000000001100011000000000000",--19804
"111110001100011000000011000000000000",--19805
"111110001110001001100011000000000000",--19806
"101111000001110001110100001000010000",--19807
"111110001110001001000011100000000000",--19808
"101111000001110010000100000101010000",--19809
"111110010000000001100011000000000000",--19810
"111110001100011000000011000000000000",--19811
"111110001110001001100011000000000000",--19812
"101111000001110001110100000111001000",--19813
"111110001110001001000011100000000000",--19814
"101111000001110010000100000100110000",--19815
"111110010000000001100011000000000000",--19816
"111110001100011000000011000000000000",--19817
"111110001110001001100011000000000000",--19818
"101111000001110001110100000110000000",--19819
"111110001110001001000011100000000000",--19820
"101111000001110010000100000100010000",--19821
"111110010000000001100011000000000000",--19822
"111110001100011000000011000000000000",--19823
"111110001110001001100011000000000000",--19824
"101111000001110001110100000100010000",--19825
"111110001110001001000011100000000000",--19826
"101111000001110010000100000011100000",--19827
"111110010000000001100011000000000000",--19828
"111110001100011000000011000000000000",--19829
"111110001110001001100011000000000000",--19830
"101111000001110010000100000010000000",--19831
"111110010000001001000100000000000000",--19832
"101111000001110010010100000010100000",--19833
"111110010010000001100011000000000000",--19834
"111110001100011000000011000000000000",--19835
"111110010000001001100011000000000000",--19836
"001001111100000001001111111111110111",--19837
"001011111100000000111111111111110110",--19838
"101110001101111000000010100000000000",--19839
"101110000011111000000001100000000000",--19840
"001001111100000111111111111111110101",--19841
"101001111100010111100000000000001100",--19842
"000111000000000000000000001101001100",--19843
"101001111100000111100000000000001100",--19844
"001101111100000111111111111111110101",--19845
"111110000110000000010001100000000000",--19846
"111110000110011000000001100000000000",--19847
"001111111100000001001111111111110110",--19848
"111110001000001000110001100000000000",--19849
"001101111100000000011111111111110111",--19850
"010100000011000000000000000000000100",--19851
"101111001001110001000011111111001001",--19852
"101111001001100001000000111111011010",--19853
"111110001000010000110001100000000000",--19854
"000101000000000000000100110110010100",--19855
"011000000011000000000000000000000011",--19856
"101111001001110001001011111111001001",--19857
"101111001001100001000000111111011010",--19858
"111110001000010000110001100000000000",--19859
"101111000001110001000100000111110000",--19860
"111110000110001001000001100000000000",--19861
"101111001001110001000011111010100010",--19862
"101111001001100001001111100110000010",--19863
"111110000110001001000001100000000000",--19864
"101110000110110000000010000000000000",--19865
"111110000110010001000001100000000000",--19866
"001111111100000001001111111111111000",--19867
"101110001001111000000010100000000001",--19868
"101111001101110001100011100011010001",--19869
"101111001101100001101011011100010111",--19870
"001011111100000000111111111111110111",--19871
"010110001101000001010000000000000010",--19872
"101111000001110000110100000101110000",--19873
"000101000000000000000100111000001111",--19874
"001111000000000001010000000100101011",--19875
"001101111100000000011111111111111001",--19876
"001111000010000001100000000000000001",--19877
"111110001010010001100010100000000000",--19878
"001101111100000000011111111111111010",--19879
"001111000010000001100000000000000001",--19880
"111110001100100000000011000000000000",--19881
"111110001010001001100010100000000000",--19882
"111110001000011000000010000000000000",--19883
"111110001010001001000010000000000001",--19884
"010110001001000000010000000000000010",--19885
"101001000000000000010000000000000001",--19886
"000101000000000000000100110110110101",--19887
"011010001001000000100000000000000010",--19888
"101001000000000000011111111111111111",--19889
"000101000000000000000100110110110101",--19890
"101000000001111000000000100000000000",--19891
"000101000000000000000100110110110110",--19892
"111110001000011000000010000000000000",--19893
"111110001000001001000010100000000000",--19894
"101111000001110001100100001011110010",--19895
"111110001100001001010011000000000000",--19896
"101111001111110001110011110100110010",--19897
"101111001111100001110001011001000011",--19898
"111110001100001001110011000000000000",--19899
"101111000001110001110100001011001000",--19900
"111110001110001001010011100000000000",--19901
"101111000001110010000100000110101000",--19902
"111110010000000001100011000000000000",--19903
"111110001100011000000011000000000000",--19904
"111110001110001001100011000000000000",--19905
"101111000001110001110100001010100010",--19906
"111110001110001001010011100000000000",--19907
"101111000001110010000100000110011000",--19908
"111110010000000001100011000000000000",--19909
"111110001100011000000011000000000000",--19910
"111110001110001001100011000000000000",--19911
"101111000001110001110100001010000000",--19912
"111110001110001001010011100000000000",--19913
"101111000001110010000100000110001000",--19914
"111110010000000001100011000000000000",--19915
"111110001100011000000011000000000000",--19916
"111110001110001001100011000000000000",--19917
"101111000001110001110100001001000100",--19918
"111110001110001001010011100000000000",--19919
"101111000001110010000100000101110000",--19920
"111110010000000001100011000000000000",--19921
"111110001100011000000011000000000000",--19922
"111110001110001001100011000000000000",--19923
"101111000001110001110100001000010000",--19924
"111110001110001001010011100000000000",--19925
"101111000001110010000100000101010000",--19926
"111110010000000001100011000000000000",--19927
"111110001100011000000011000000000000",--19928
"111110001110001001100011000000000000",--19929
"101111000001110001110100000111001000",--19930
"111110001110001001010011100000000000",--19931
"101111000001110010000100000100110000",--19932
"111110010000000001100011000000000000",--19933
"111110001100011000000011000000000000",--19934
"111110001110001001100011000000000000",--19935
"101111000001110001110100000110000000",--19936
"111110001110001001010011100000000000",--19937
"101111000001110010000100000100010000",--19938
"111110010000000001100011000000000000",--19939
"111110001100011000000011000000000000",--19940
"111110001110001001100011000000000000",--19941
"101111000001110001110100000100010000",--19942
"111110001110001001010011100000000000",--19943
"101111000001110010000100000011100000",--19944
"111110010000000001100011000000000000",--19945
"111110001100011000000011000000000000",--19946
"111110001110001001100011000000000000",--19947
"101111000001110010000100000010000000",--19948
"111110010000001001010100000000000000",--19949
"101111000001110010010100000010100000",--19950
"111110010010000001100011000000000000",--19951
"111110001100011000000011000000000000",--19952
"111110010000001001100011000000000000",--19953
"001001111100000000011111111111110110",--19954
"001011111100000001001111111111110101",--19955
"101110001011111000000010000000000000",--19956
"101110000011111000000001100000000000",--19957
"101110001101111000000010100000000000",--19958
"001001111100000111111111111111110100",--19959
"101001111100010111100000000000001101",--19960
"000111000000000000000000001101001100",--19961
"101001111100000111100000000000001101",--19962
"001101111100000111111111111111110100",--19963
"111110000110000000010001100000000000",--19964
"111110000110011000000001100000000000",--19965
"001111111100000001001111111111110101",--19966
"111110001000001000110001100000000000",--19967
"001101111100000000011111111111110110",--19968
"010100000011000000000000000000000100",--19969
"101111001001110001000011111111001001",--19970
"101111001001100001000000111111011010",--19971
"111110001000010000110001100000000000",--19972
"000101000000000000000100111000001010",--19973
"011000000011000000000000000000000011",--19974
"101111001001110001001011111111001001",--19975
"101111001001100001000000111111011010",--19976
"111110001000010000110001100000000000",--19977
"101111000001110001000100000111110000",--19978
"111110000110001001000001100000000000",--19979
"101111001001110001000011111010100010",--19980
"101111001001100001001111100110000010",--19981
"111110000110001001000001100000000000",--19982
"101110000110110000000010000000000000",--19983
"111110000110010001000001100000000000",--19984
"101111001001110001000011111000011001",--19985
"101111001001100001001001100110011010",--19986
"101111000001110001010011111100000000",--19987
"001111111100000001101111111111110111",--19988
"111110001010010001100010100000000000",--19989
"111110001010001001010010100000000000",--19990
"111110001000010001010010000000000000",--19991
"101111000001110001010011111100000000",--19992
"111110001010010000110001100000000000",--19993
"111110000110001000110001100000000000",--19994
"111110001000010000110001100000000000",--19995
"011010000111000000000000000000000001",--19996
"101110000001111000000001100000000000",--19997
"101111000001110001000100001101111111",--19998
"111110001000001000110001100000000000",--19999
"101111001001110001000100000001010101",--20000
"101111001001100001000101010101010101",--20001
"111110000110001001000001100000000000",--20002
"001011000000000000110000000100100101",--20003
"001101000000000000100000000100110000",--20004
"001101000100000000010000000000000000",--20005
"001101000010000000110000000000000000",--20006
"010011000111000000000000000010110100",--20007
"001001111100000000011111111111111010",--20008
"001001111100000000101111111111111001",--20009
"010011000111011000110000000010100010",--20010
"001101000110000001000000000101101101",--20011
"001111000000000000110000000100101010",--20012
"001101001000000001010000000000000101",--20013
"001111001010000001000000000000000000",--20014
"111110000110010001000001100000000000",--20015
"001111000000000001000000000100101011",--20016
"001111001010000001010000000000000001",--20017
"111110001000010001010010000000000000",--20018
"001111000000000001010000000100101100",--20019
"001111001010000001100000000000000010",--20020
"111110001010010001100010100000000000",--20021
"001101000110000000110000000010111110",--20022
"001101001000000001010000000000000001",--20023
"011111001011000000010000000000110111",--20024
"001111000110000001100000000000000000",--20025
"111110001100010000110011000000000000",--20026
"001111000110000001110000000000000001",--20027
"111110001100001001110011000000000000",--20028
"001111000000000001110000000011111011",--20029
"111110001100001001110011100000000000",--20030
"111110001110000001000011100000000001",--20031
"001101001000000001000000000000000100",--20032
"001111001000000010000000000000000001",--20033
"010110010001000001110000000000000111",--20034
"001111000000000001110000000011111100",--20035
"111110001100001001110011100000000000",--20036
"111110001110000001010011100000000001",--20037
"001111001000000010000000000000000010",--20038
"010110010001000001110000000000000010",--20039
"001111000110000001110000000000000001",--20040
"011110001111000000000000000000100100",--20041
"001111000110000001100000000000000010",--20042
"111110001100010001000011000000000000",--20043
"001111000110000001110000000000000011",--20044
"111110001100001001110011000000000000",--20045
"001111000000000001110000000011111010",--20046
"111110001100001001110011100000000000",--20047
"111110001110000000110011100000000001",--20048
"001111001000000010000000000000000000",--20049
"010110010001000001110000000000000111",--20050
"001111000000000001110000000011111100",--20051
"111110001100001001110011100000000000",--20052
"111110001110000001010011100000000001",--20053
"001111001000000010000000000000000010",--20054
"010110010001000001110000000000000010",--20055
"001111000110000001110000000000000011",--20056
"011110001111000000000000000000010010",--20057
"001111000110000001100000000000000100",--20058
"111110001100010001010010100000000000",--20059
"001111000110000001100000000000000101",--20060
"111110001010001001100010100000000000",--20061
"001111000000000001100000000011111010",--20062
"111110001010001001100011000000000000",--20063
"111110001100000000110001100000000001",--20064
"001111001000000001100000000000000000",--20065
"010110001101000000110000000001100001",--20066
"001111000000000000110000000011111011",--20067
"111110001010001000110001100000000000",--20068
"111110000110000001000001100000000001",--20069
"001111001000000001000000000000000001",--20070
"010110001001000000110000000001011100",--20071
"001111000110000000110000000000000101",--20072
"010010000111000000000000000001011010",--20073
"001011000000000001010000000100101111",--20074
"000101000000000000000100111010111000",--20075
"001011000000000001100000000100101111",--20076
"000101000000000000000100111010111000",--20077
"001011000000000001100000000100101111",--20078
"000101000000000000000100111010111000",--20079
"011111001011000000100000000000001100",--20080
"001111000110000001100000000000000000",--20081
"011010001101000000000000000001010001",--20082
"001111000110000001100000000000000001",--20083
"111110001100001000110001100000000000",--20084
"001111000110000001100000000000000010",--20085
"111110001100001001000010000000000000",--20086
"111110000110000001000001100000000000",--20087
"001111000110000001000000000000000011",--20088
"111110001000001001010010000000000000",--20089
"111110000110000001000001100000000000",--20090
"001011000000000000110000000100101111",--20091
"000101000000000000000100111010111000",--20092
"001111000110000001100000000000000000",--20093
"010010001101000000000000000001000101",--20094
"001111000110000001110000000000000001",--20095
"111110001110001000110011100000000000",--20096
"001111000110000010000000000000000010",--20097
"111110010000001001000100000000000000",--20098
"111110001110000010000011100000000000",--20099
"001111000110000010000000000000000011",--20100
"111110010000001001010100000000000000",--20101
"111110001110000010000011100000000000",--20102
"111110000110001000110100000000000000",--20103
"001101001000000001100000000000000100",--20104
"001111001100000010010000000000000000",--20105
"111110010000001010010100000000000000",--20106
"111110001000001001000100100000000000",--20107
"001111001100000010100000000000000001",--20108
"111110010010001010100100100000000000",--20109
"111110010000000010010100000000000000",--20110
"111110001010001001010100100000000000",--20111
"001111001100000010100000000000000010",--20112
"111110010010001010100100100000000000",--20113
"111110010000000010010100000000000000",--20114
"001101001000000001100000000000000011",--20115
"011100001101000000000000000000000011",--20116
"101110010001111000000001100000000000",--20117
"011111001011000000110000000000010000",--20118
"000101000000000000000100111010100110",--20119
"111110001000001001010100100000000000",--20120
"001101001000000001100000000000001001",--20121
"001111001100000010100000000000000000",--20122
"111110010010001010100100100000000000",--20123
"111110010000000010010100000000000000",--20124
"111110001010001000110010100000000000",--20125
"001111001100000010010000000000000001",--20126
"111110001010001010010010100000000000",--20127
"111110010000000001010010100000000000",--20128
"111110000110001001000001100000000000",--20129
"001111001100000001000000000000000010",--20130
"111110000110001001000001100000000000",--20131
"111110001010000000110001100000000000",--20132
"011111001011000000110000000000000001",--20133
"111110000110010000010001100000000000",--20134
"111110001110001001110010000000000000",--20135
"111110001100001000110001100000000000",--20136
"111110001000010000110001100000000000",--20137
"010110000111000000000000000000011001",--20138
"001101001000000001000000000000000110",--20139
"011100001001000000000000000000000110",--20140
"111110000110100000000001100000000000",--20141
"111110001110010000110001100000000000",--20142
"001111000110000001000000000000000100",--20143
"111110000110001001000001100000000000",--20144
"001011000000000000110000000100101111",--20145
"000101000000000000000100111010111000",--20146
"111110000110100000000001100000000000",--20147
"111110001110000000110001100000000000",--20148
"001111000110000001000000000000000100",--20149
"111110000110001001000001100000000000",--20150
"001011000000000000110000000100101111",--20151
"001111000000000000110000000100101111",--20152
"101111001001110001001011110111001100",--20153
"101111001001100001001100110011001101",--20154
"010110001001000000110000000000001000",--20155
"101000000011111000000001000000000000",--20156
"101001000000000000010000000000000001",--20157
"001001111100000111111111111111111000",--20158
"101001111100010111100000000000001001",--20159
"000111000000000000000000110101111110",--20160
"101001111100000111100000000000001001",--20161
"001101111100000111111111111111111000",--20162
"011100000011000000000000000000001001",--20163
"101001000000000000010000000000000001",--20164
"001101111100000000101111111111111001",--20165
"001001111100000111111111111111111000",--20166
"101001111100010111100000000000001001",--20167
"000111000000000000000000111111111011",--20168
"101001111100000111100000000000001001",--20169
"001101111100000111111111111111111000",--20170
"011100000011000000000000001011111100",--20171
"000101000000000000000100111011011100",--20172
"101001000000000000010000000000000001",--20173
"001101111100000000101111111111111010",--20174
"001001111100000111111111111111111000",--20175
"101001111100010111100000000000001001",--20176
"000111000000000000000000110101111110",--20177
"101001111100000111100000000000001001",--20178
"001101111100000111111111111111111000",--20179
"011100000011000000000000001011110011",--20180
"101001000000000000010000000000000001",--20181
"001101111100000000101111111111111001",--20182
"101001111100010111100000000000001001",--20183
"000111000000000000000000111111111011",--20184
"101001111100000111100000000000001001",--20185
"001101111100000111111111111111111000",--20186
"011100000011000000000000001011101100",--20187
"101111000111110000111011101111011010",--20188
"101111000111100000110111010000001101",--20189
"001111111100000001001111111111111101",--20190
"111110001000001000110001100000000000",--20191
"001111000000000001000000000100100110",--20192
"001111000000000001010000000101100100",--20193
"111110001000001001010010000000000000",--20194
"001111000000000001010000000100100111",--20195
"001111000000000001100000000101100101",--20196
"111110001010001001100010100000000000",--20197
"111110001000000001010010000000000000",--20198
"001111000000000001010000000100101000",--20199
"001111000000000001100000000101100110",--20200
"111110001010001001100010100000000000",--20201
"111110001000000001010010000000000010",--20202
"010110001001000000000000000000000001",--20203
"000101000000000000000100111011101110",--20204
"101110000001111000000010000000000000",--20205
"111110000110001001000001100000000000",--20206
"001101111100000000011111111111111011",--20207
"001101000010000000010000000000000111",--20208
"001111000010000001000000000000000000",--20209
"111110000110001001000001100000000000",--20210
"001111000000000001000000000100100000",--20211
"001111000000000001010000000100100011",--20212
"111110000110001001010010100000000000",--20213
"111110001000000001010010000000000000",--20214
"001011000000000001000000000100100000",--20215
"001111000000000001000000000100100001",--20216
"001111000000000001010000000100100100",--20217
"111110000110001001010010100000000000",--20218
"111110001000000001010010000000000000",--20219
"001011000000000001000000000100100001",--20220
"001111000000000001000000000100100010",--20221
"001111000000000001010000000100100101",--20222
"111110000110001001010001100000000000",--20223
"111110001000000000110001100000000000",--20224
"001011000000000000110000000100100010",--20225
"000101000000000000000101000111001000",--20226
"001101000010000000110000000001110110",--20227
"101111001001110001000100111001101110",--20228
"101111001001100001000110101100101000",--20229
"001011000000000001000000000100101101",--20230
"001101000000000000100000000100110000",--20231
"001011111100000000111111111111111101",--20232
"001001111100000000111111111111111100",--20233
"101000000001111000000000100000000000",--20234
"001001111100000111111111111111111011",--20235
"101001111100010111100000000000000110",--20236
"000111000000000000000010110111111111",--20237
"101001111100000111100000000000000110",--20238
"001101111100000111111111111111111011",--20239
"001111000000000000110000000100101101",--20240
"101111001001110001001011110111001100",--20241
"101111001001100001001100110011001101",--20242
"010110000111000001000000001010110100",--20243
"101111001001110001000100110010111110",--20244
"101111001001100001001011110000100000",--20245
"010110001001000000110000001010110001",--20246
"001101000000000000010000000100101001",--20247
"001101000010000000010000000101101101",--20248
"001101000010000000100000000000000001",--20249
"011111000101000000010000000000010011",--20250
"001101111100000000101111111111111100",--20251
"001101000100000000100000000000000000",--20252
"001101000000000000110000000100101110",--20253
"001011000000000000000000000100100110",--20254
"001011000000000000000000000100100111",--20255
"001011000000000000000000000100101000",--20256
"101001000110010001000000000000000001",--20257
"101001000110010000110000000000000001",--20258
"001110000100000000110001100000000000",--20259
"011110000111000000000000000000000010",--20260
"101110000001111000000001100000000000",--20261
"000101000000000000000100111100101011",--20262
"010110000111000000000000000000000010",--20263
"101110000011111000000001100000000000",--20264
"000101000000000000000100111100101011",--20265
"101110000101111000000001100000000000",--20266
"101110000111111000000001100000000010",--20267
"001011001000000000110000000100100110",--20268
"000101000000000000000100111110000100",--20269
"011111000101000000100000000000001000",--20270
"001101000010000000100000000000000100",--20271
"001111000100010000110000000000000000",--20272
"001011000000000000110000000100100110",--20273
"001111000100010000110000000000000001",--20274
"001011000000000000110000000100100111",--20275
"001111000100010000110000000000000010",--20276
"001011000000000000110000000100101000",--20277
"000101000000000000000100111110000100",--20278
"001111000000000000110000000100101010",--20279
"001101000010000000100000000000000101",--20280
"001111000100000001000000000000000000",--20281
"111110000110010001000001100000000000",--20282
"001111000000000001000000000100101011",--20283
"001111000100000001010000000000000001",--20284
"111110001000010001010010000000000000",--20285
"001111000000000001010000000100101100",--20286
"001111000100000001100000000000000010",--20287
"111110001010010001100010100000000000",--20288
"001101000010000000100000000000000100",--20289
"001111000100000001100000000000000000",--20290
"111110000110001001100011000000000000",--20291
"001111000100000001110000000000000001",--20292
"111110001000001001110011100000000000",--20293
"001111000100000010000000000000000010",--20294
"111110001010001010000100000000000000",--20295
"001101000010000000100000000000000011",--20296
"011100000101000000000000000000000100",--20297
"001011000000000001100000000100100110",--20298
"001011000000000001110000000100100111",--20299
"001011000000000010000000000100101000",--20300
"000101000000000000000100111101101010",--20301
"001101000010000000100000000000001001",--20302
"001111000100000010010000000000000010",--20303
"111110001000001010010100100000000000",--20304
"001111000100000010100000000000000001",--20305
"111110001010001010100101000000000000",--20306
"111110010010000010100100100000000000",--20307
"101111000001110010100011111100000000",--20308
"111110010010001010100100100000000000",--20309
"111110001100000010010011000000000000",--20310
"001011000000000001100000000100100110",--20311
"001111000100000001100000000000000010",--20312
"111110000110001001100011000000000000",--20313
"001111000100000010010000000000000000",--20314
"111110001010001010010010100000000000",--20315
"111110001100000001010010100000000000",--20316
"101111000001110001100011111100000000",--20317
"111110001010001001100010100000000000",--20318
"111110001110000001010010100000000000",--20319
"001011000000000001010000000100100111",--20320
"001111000100000001010000000000000001",--20321
"111110000110001001010001100000000000",--20322
"001111000100000001010000000000000000",--20323
"111110001000001001010010000000000000",--20324
"111110000110000001000001100000000000",--20325
"101111000001110001000011111100000000",--20326
"111110000110001001000001100000000000",--20327
"111110010000000000110001100000000000",--20328
"001011000000000000110000000100101000",--20329
"001111000000000000110000000100100110",--20330
"111110000110001000110001100000000000",--20331
"001111000000000001000000000100100111",--20332
"111110001000001001000010000000000000",--20333
"111110000110000001000001100000000000",--20334
"001111000000000001000000000100101000",--20335
"111110001000001001000010000000000000",--20336
"111110000110000001000001100000000000",--20337
"111110000110100000000001100000000000",--20338
"011110000111000000000000000000000010",--20339
"101110000011111000000001100000000000",--20340
"000101000000000000000100111101111011",--20341
"001101000010000000100000000000000110",--20342
"011100000101000000000000000000000010",--20343
"111110000110011000000001100000000000",--20344
"000101000000000000000100111101111011",--20345
"111110000110011000000001100000000010",--20346
"001111000000000001000000000100100110",--20347
"111110001000001000110010000000000000",--20348
"001011000000000001000000000100100110",--20349
"001111000000000001000000000100100111",--20350
"111110001000001000110010000000000000",--20351
"001011000000000001000000000100100111",--20352
"001111000000000001000000000100101000",--20353
"111110001000001000110001100000000000",--20354
"001011000000000000110000000100101000",--20355
"001101000010000000100000000000000000",--20356
"001101000010000000110000000000001000",--20357
"001111000110000000110000000000000000",--20358
"001011000000000000110000000100100011",--20359
"001111000110000000110000000000000001",--20360
"001011000000000000110000000100100100",--20361
"001111000110000000110000000000000010",--20362
"001011000000000000110000000100100101",--20363
"001001111100000000011111111111111011",--20364
"011111000101000000010000000000100011",--20365
"001111000000000000110000000100101010",--20366
"001101000010000000100000000000000101",--20367
"001111000100000001000000000000000000",--20368
"111110000110010001000001100000000000",--20369
"101111001001110001000011110101001100",--20370
"101111001001100001001100110011001101",--20371
"111110000110001001000010000000000000",--20372
"101110001000110000000010000000000000",--20373
"101111000001110001010100000110100000",--20374
"111110001000001001010010000000000000",--20375
"111110000110010001000001100000000000",--20376
"101111000001110001000100000100100000",--20377
"001111000000000001010000000100101100",--20378
"001111000100000001100000000000000010",--20379
"111110001010010001100010100000000000",--20380
"101111001101110001100011110101001100",--20381
"101111001101100001101100110011001101",--20382
"111110001010001001100011000000000000",--20383
"101110001100110000000011000000000000",--20384
"101111000001110001110100000110100000",--20385
"111110001100001001110011000000000000",--20386
"111110001010010001100010100000000000",--20387
"101111000001110001100100000100100000",--20388
"010110001001000000110000000000000101",--20389
"010110001101000001010000000000000010",--20390
"101111000001110000110100001101111111",--20391
"000101000000000000000100111110101111",--20392
"101110000001111000000001100000000000",--20393
"000101000000000000000100111110101111",--20394
"010110001101000001010000000000000010",--20395
"101110000001111000000001100000000000",--20396
"000101000000000000000100111110101111",--20397
"101111000001110000110100001101111111",--20398
"001011000000000000110000000100100100",--20399
"000101000000000000000101000011101010",--20400
"011111000101000000100000000000001111",--20401
"001111000000000000110000000100101011",--20402
"101111000001110001000011111010000000",--20403
"111110000110001001000001100000000000",--20404
"001001111100000111111111111111111010",--20405
"000111000000000000000111011000000010",--20406
"001101111100000111111111111111111010",--20407
"111110000110001000110001100000000000",--20408
"101111000001110001000100001101111111",--20409
"111110001000001000110010000000000000",--20410
"001011000000000001000000000100100011",--20411
"101111000001110001000100001101111111",--20412
"111110000110010000010001100000000010",--20413
"111110001000001000110001100000000000",--20414
"001011000000000000110000000100100100",--20415
"000101000000000000000101000011101010",--20416
"011111000101000000110000000000011111",--20417
"001111000000000000110000000100101010",--20418
"001101000010000000100000000000000101",--20419
"001111000100000001000000000000000000",--20420
"111110000110010001000001100000000000",--20421
"001111000000000001000000000100101100",--20422
"001111000100000001010000000000000010",--20423
"111110001000010001010010000000000000",--20424
"111110000110001000110001100000000000",--20425
"111110001000001001000010000000000000",--20426
"111110000110000001000001100000000000",--20427
"111110000110100000000001100000000000",--20428
"101111001001110001000011110111001100",--20429
"101111001001100001001100110011001100",--20430
"111110000110001001000001100000000000",--20431
"101110000110110000000010000000000000",--20432
"111110000110010001000001100000000000",--20433
"101111001001110001000100000001001001",--20434
"101111001001100001000000111111011011",--20435
"111110000110001001000001100000000000",--20436
"001001111100000111111111111111111010",--20437
"000111000000000000000111010110111000",--20438
"001101111100000111111111111111111010",--20439
"111110000110001000110001100000000000",--20440
"101111000001110001000100001101111111",--20441
"111110000110001001000010000000000000",--20442
"001011000000000001000000000100100100",--20443
"111110000110010000010001100000000010",--20444
"101111000001110001000100001101111111",--20445
"111110000110001001000001100000000000",--20446
"001011000000000000110000000100100101",--20447
"000101000000000000000101000011101010",--20448
"011111000101000001000000000100001000",--20449
"001111000000000000110000000100101010",--20450
"001101000010000000100000000000000101",--20451
"001111000100000001000000000000000000",--20452
"111110000110010001000001100000000000",--20453
"001101000010000000110000000000000100",--20454
"001111000110000001000000000000000000",--20455
"111110001000100000000010000000000000",--20456
"111110000110001001000001100000000000",--20457
"001111000000000001000000000100101100",--20458
"001111000100000001010000000000000010",--20459
"111110001000010001010010000000000000",--20460
"001111000110000001010000000000000010",--20461
"111110001010100000000010100000000000",--20462
"111110001000001001010010000000000000",--20463
"111110000110001000110010100000000000",--20464
"111110001000001001000011000000000000",--20465
"111110001010000001100010100000000000",--20466
"101110000111111000000011000000000001",--20467
"101111001111110001110011100011010001",--20468
"101111001111100001111011011100010111",--20469
"001001111100000000111111111111111010",--20470
"001001111100000000101111111111111001",--20471
"001011111100000001011111111111111000",--20472
"010110001111000001100000000000000010",--20473
"101111000001110000110100000101110000",--20474
"000101000000000000000101000001011111",--20475
"111110000110011000000001100000000000",--20476
"111110001000001000110001100000000001",--20477
"010110000111000000010000000000000010",--20478
"101001000000000001000000000000000001",--20479
"000101000000000000000101000000000110",--20480
"011010000111000000100000000000000010",--20481
"101001000000000001001111111111111111",--20482
"000101000000000000000101000000000110",--20483
"101000000001111000000010000000000000",--20484
"000101000000000000000101000000000111",--20485
"111110000110011000000001100000000000",--20486
"111110000110001000110010000000000000",--20487
"101111000001110001100100001011110010",--20488
"111110001100001001000011000000000000",--20489
"101111001111110001110011110100110010",--20490
"101111001111100001110001011001000011",--20491
"111110001100001001110011000000000000",--20492
"101111000001110001110100001011001000",--20493
"111110001110001001000011100000000000",--20494
"101111000001110010000100000110101000",--20495
"111110010000000001100011000000000000",--20496
"111110001100011000000011000000000000",--20497
"111110001110001001100011000000000000",--20498
"101111000001110001110100001010100010",--20499
"111110001110001001000011100000000000",--20500
"101111000001110010000100000110011000",--20501
"111110010000000001100011000000000000",--20502
"111110001100011000000011000000000000",--20503
"111110001110001001100011000000000000",--20504
"101111000001110001110100001010000000",--20505
"111110001110001001000011100000000000",--20506
"101111000001110010000100000110001000",--20507
"111110010000000001100011000000000000",--20508
"111110001100011000000011000000000000",--20509
"111110001110001001100011000000000000",--20510
"101111000001110001110100001001000100",--20511
"111110001110001001000011100000000000",--20512
"101111000001110010000100000101110000",--20513
"111110010000000001100011000000000000",--20514
"111110001100011000000011000000000000",--20515
"111110001110001001100011000000000000",--20516
"101111000001110001110100001000010000",--20517
"111110001110001001000011100000000000",--20518
"101111000001110010000100000101010000",--20519
"111110010000000001100011000000000000",--20520
"111110001100011000000011000000000000",--20521
"111110001110001001100011000000000000",--20522
"101111000001110001110100000111001000",--20523
"111110001110001001000011100000000000",--20524
"101111000001110010000100000100110000",--20525
"111110010000000001100011000000000000",--20526
"111110001100011000000011000000000000",--20527
"111110001110001001100011000000000000",--20528
"101111000001110001110100000110000000",--20529
"111110001110001001000011100000000000",--20530
"101111000001110010000100000100010000",--20531
"111110010000000001100011000000000000",--20532
"111110001100011000000011000000000000",--20533
"111110001110001001100011000000000000",--20534
"101111000001110001110100000100010000",--20535
"111110001110001001000011100000000000",--20536
"101111000001110010000100000011100000",--20537
"111110010000000001100011000000000000",--20538
"111110001100011000000011000000000000",--20539
"111110001110001001100011000000000000",--20540
"101111000001110010000100000010000000",--20541
"111110010000001001000100000000000000",--20542
"101111000001110010010100000010100000",--20543
"111110010010000001100011000000000000",--20544
"111110001100011000000011000000000000",--20545
"111110010000001001100011000000000000",--20546
"001001111100000001001111111111110111",--20547
"001011111100000000111111111111110110",--20548
"101110001101111000000010100000000000",--20549
"101110000011111000000001100000000000",--20550
"001001111100000111111111111111110101",--20551
"101001111100010111100000000000001100",--20552
"000111000000000000000000001101001100",--20553
"101001111100000111100000000000001100",--20554
"001101111100000111111111111111110101",--20555
"111110000110000000010001100000000000",--20556
"111110000110011000000001100000000000",--20557
"001111111100000001001111111111110110",--20558
"111110001000001000110001100000000000",--20559
"001101111100000000011111111111110111",--20560
"010100000011000000000000000000000100",--20561
"101111001001110001000011111111001001",--20562
"101111001001100001000000111111011010",--20563
"111110001000010000110001100000000000",--20564
"000101000000000000000101000001011010",--20565
"011000000011000000000000000000000011",--20566
"101111001001110001001011111111001001",--20567
"101111001001100001000000111111011010",--20568
"111110001000010000110001100000000000",--20569
"101111000001110001000100000111110000",--20570
"111110000110001001000001100000000000",--20571
"101111001001110001000011111010100010",--20572
"101111001001100001001111100110000010",--20573
"111110000110001001000001100000000000",--20574
"101110000110110000000010000000000000",--20575
"111110000110010001000001100000000000",--20576
"001111111100000001001111111111111000",--20577
"101110001001111000000010100000000001",--20578
"101111001101110001100011100011010001",--20579
"101111001101100001101011011100010111",--20580
"001011111100000000111111111111110111",--20581
"010110001101000001010000000000000010",--20582
"101111000001110000110100000101110000",--20583
"000101000000000000000101000011010101",--20584
"001111000000000001010000000100101011",--20585
"001101111100000000011111111111111001",--20586
"001111000010000001100000000000000001",--20587
"111110001010010001100010100000000000",--20588
"001101111100000000011111111111111010",--20589
"001111000010000001100000000000000001",--20590
"111110001100100000000011000000000000",--20591
"111110001010001001100010100000000000",--20592
"111110001000011000000010000000000000",--20593
"111110001010001001000010000000000001",--20594
"010110001001000000010000000000000010",--20595
"101001000000000000010000000000000001",--20596
"000101000000000000000101000001111011",--20597
"011010001001000000100000000000000010",--20598
"101001000000000000011111111111111111",--20599
"000101000000000000000101000001111011",--20600
"101000000001111000000000100000000000",--20601
"000101000000000000000101000001111100",--20602
"111110001000011000000010000000000000",--20603
"111110001000001001000010100000000000",--20604
"101111000001110001100100001011110010",--20605
"111110001100001001010011000000000000",--20606
"101111001111110001110011110100110010",--20607
"101111001111100001110001011001000011",--20608
"111110001100001001110011000000000000",--20609
"101111000001110001110100001011001000",--20610
"111110001110001001010011100000000000",--20611
"101111000001110010000100000110101000",--20612
"111110010000000001100011000000000000",--20613
"111110001100011000000011000000000000",--20614
"111110001110001001100011000000000000",--20615
"101111000001110001110100001010100010",--20616
"111110001110001001010011100000000000",--20617
"101111000001110010000100000110011000",--20618
"111110010000000001100011000000000000",--20619
"111110001100011000000011000000000000",--20620
"111110001110001001100011000000000000",--20621
"101111000001110001110100001010000000",--20622
"111110001110001001010011100000000000",--20623
"101111000001110010000100000110001000",--20624
"111110010000000001100011000000000000",--20625
"111110001100011000000011000000000000",--20626
"111110001110001001100011000000000000",--20627
"101111000001110001110100001001000100",--20628
"111110001110001001010011100000000000",--20629
"101111000001110010000100000101110000",--20630
"111110010000000001100011000000000000",--20631
"111110001100011000000011000000000000",--20632
"111110001110001001100011000000000000",--20633
"101111000001110001110100001000010000",--20634
"111110001110001001010011100000000000",--20635
"101111000001110010000100000101010000",--20636
"111110010000000001100011000000000000",--20637
"111110001100011000000011000000000000",--20638
"111110001110001001100011000000000000",--20639
"101111000001110001110100000111001000",--20640
"111110001110001001010011100000000000",--20641
"101111000001110010000100000100110000",--20642
"111110010000000001100011000000000000",--20643
"111110001100011000000011000000000000",--20644
"111110001110001001100011000000000000",--20645
"101111000001110001110100000110000000",--20646
"111110001110001001010011100000000000",--20647
"101111000001110010000100000100010000",--20648
"111110010000000001100011000000000000",--20649
"111110001100011000000011000000000000",--20650
"111110001110001001100011000000000000",--20651
"101111000001110001110100000100010000",--20652
"111110001110001001010011100000000000",--20653
"101111000001110010000100000011100000",--20654
"111110010000000001100011000000000000",--20655
"111110001100011000000011000000000000",--20656
"111110001110001001100011000000000000",--20657
"101111000001110010000100000010000000",--20658
"111110010000001001010100000000000000",--20659
"101111000001110010010100000010100000",--20660
"111110010010000001100011000000000000",--20661
"111110001100011000000011000000000000",--20662
"111110010000001001100011000000000000",--20663
"001001111100000000011111111111110110",--20664
"001011111100000001001111111111110101",--20665
"101110001011111000000010000000000000",--20666
"101110000011111000000001100000000000",--20667
"101110001101111000000010100000000000",--20668
"001001111100000111111111111111110100",--20669
"101001111100010111100000000000001101",--20670
"000111000000000000000000001101001100",--20671
"101001111100000111100000000000001101",--20672
"001101111100000111111111111111110100",--20673
"111110000110000000010001100000000000",--20674
"111110000110011000000001100000000000",--20675
"001111111100000001001111111111110101",--20676
"111110001000001000110001100000000000",--20677
"001101111100000000011111111111110110",--20678
"010100000011000000000000000000000100",--20679
"101111001001110001000011111111001001",--20680
"101111001001100001000000111111011010",--20681
"111110001000010000110001100000000000",--20682
"000101000000000000000101000011010000",--20683
"011000000011000000000000000000000011",--20684
"101111001001110001001011111111001001",--20685
"101111001001100001000000111111011010",--20686
"111110001000010000110001100000000000",--20687
"101111000001110001000100000111110000",--20688
"111110000110001001000001100000000000",--20689
"101111001001110001000011111010100010",--20690
"101111001001100001001111100110000010",--20691
"111110000110001001000001100000000000",--20692
"101110000110110000000010000000000000",--20693
"111110000110010001000001100000000000",--20694
"101111001001110001000011111000011001",--20695
"101111001001100001001001100110011010",--20696
"101111000001110001010011111100000000",--20697
"001111111100000001101111111111110111",--20698
"111110001010010001100010100000000000",--20699
"111110001010001001010010100000000000",--20700
"111110001000010001010010000000000000",--20701
"101111000001110001010011111100000000",--20702
"111110001010010000110001100000000000",--20703
"111110000110001000110001100000000000",--20704
"111110001000010000110001100000000000",--20705
"011010000111000000000000000000000001",--20706
"101110000001111000000001100000000000",--20707
"101111000001110001000100001101111111",--20708
"111110001000001000110001100000000000",--20709
"101111001001110001000100000001010101",--20710
"101111001001100001000101010101010101",--20711
"111110000110001001000001100000000000",--20712
"001011000000000000110000000100100101",--20713
"001101000000000000100000000100110000",--20714
"001101000100000000010000000000000000",--20715
"001101000010000000110000000000000000",--20716
"010011000111000000000000000010110100",--20717
"001001111100000000011111111111111010",--20718
"001001111100000000101111111111111001",--20719
"010011000111011000110000000010100010",--20720
"001101000110000001000000000101101101",--20721
"001111000000000000110000000100101010",--20722
"001101001000000001010000000000000101",--20723
"001111001010000001000000000000000000",--20724
"111110000110010001000001100000000000",--20725
"001111000000000001000000000100101011",--20726
"001111001010000001010000000000000001",--20727
"111110001000010001010010000000000000",--20728
"001111000000000001010000000100101100",--20729
"001111001010000001100000000000000010",--20730
"111110001010010001100010100000000000",--20731
"001101000110000000110000000010111110",--20732
"001101001000000001010000000000000001",--20733
"011111001011000000010000000000110111",--20734
"001111000110000001100000000000000000",--20735
"111110001100010000110011000000000000",--20736
"001111000110000001110000000000000001",--20737
"111110001100001001110011000000000000",--20738
"001111000000000001110000000011111011",--20739
"111110001100001001110011100000000000",--20740
"111110001110000001000011100000000001",--20741
"001101001000000001000000000000000100",--20742
"001111001000000010000000000000000001",--20743
"010110010001000001110000000000000111",--20744
"001111000000000001110000000011111100",--20745
"111110001100001001110011100000000000",--20746
"111110001110000001010011100000000001",--20747
"001111001000000010000000000000000010",--20748
"010110010001000001110000000000000010",--20749
"001111000110000001110000000000000001",--20750
"011110001111000000000000000000100100",--20751
"001111000110000001100000000000000010",--20752
"111110001100010001000011000000000000",--20753
"001111000110000001110000000000000011",--20754
"111110001100001001110011000000000000",--20755
"001111000000000001110000000011111010",--20756
"111110001100001001110011100000000000",--20757
"111110001110000000110011100000000001",--20758
"001111001000000010000000000000000000",--20759
"010110010001000001110000000000000111",--20760
"001111000000000001110000000011111100",--20761
"111110001100001001110011100000000000",--20762
"111110001110000001010011100000000001",--20763
"001111001000000010000000000000000010",--20764
"010110010001000001110000000000000010",--20765
"001111000110000001110000000000000011",--20766
"011110001111000000000000000000010010",--20767
"001111000110000001100000000000000100",--20768
"111110001100010001010010100000000000",--20769
"001111000110000001100000000000000101",--20770
"111110001010001001100010100000000000",--20771
"001111000000000001100000000011111010",--20772
"111110001010001001100011000000000000",--20773
"111110001100000000110001100000000001",--20774
"001111001000000001100000000000000000",--20775
"010110001101000000110000000001100001",--20776
"001111000000000000110000000011111011",--20777
"111110001010001000110001100000000000",--20778
"111110000110000001000001100000000001",--20779
"001111001000000001000000000000000001",--20780
"010110001001000000110000000001011100",--20781
"001111000110000000110000000000000101",--20782
"010010000111000000000000000001011010",--20783
"001011000000000001010000000100101111",--20784
"000101000000000000000101000101111110",--20785
"001011000000000001100000000100101111",--20786
"000101000000000000000101000101111110",--20787
"001011000000000001100000000100101111",--20788
"000101000000000000000101000101111110",--20789
"011111001011000000100000000000001100",--20790
"001111000110000001100000000000000000",--20791
"011010001101000000000000000001010001",--20792
"001111000110000001100000000000000001",--20793
"111110001100001000110001100000000000",--20794
"001111000110000001100000000000000010",--20795
"111110001100001001000010000000000000",--20796
"111110000110000001000001100000000000",--20797
"001111000110000001000000000000000011",--20798
"111110001000001001010010000000000000",--20799
"111110000110000001000001100000000000",--20800
"001011000000000000110000000100101111",--20801
"000101000000000000000101000101111110",--20802
"001111000110000001100000000000000000",--20803
"010010001101000000000000000001000101",--20804
"001111000110000001110000000000000001",--20805
"111110001110001000110011100000000000",--20806
"001111000110000010000000000000000010",--20807
"111110010000001001000100000000000000",--20808
"111110001110000010000011100000000000",--20809
"001111000110000010000000000000000011",--20810
"111110010000001001010100000000000000",--20811
"111110001110000010000011100000000000",--20812
"111110000110001000110100000000000000",--20813
"001101001000000001100000000000000100",--20814
"001111001100000010010000000000000000",--20815
"111110010000001010010100000000000000",--20816
"111110001000001001000100100000000000",--20817
"001111001100000010100000000000000001",--20818
"111110010010001010100100100000000000",--20819
"111110010000000010010100000000000000",--20820
"111110001010001001010100100000000000",--20821
"001111001100000010100000000000000010",--20822
"111110010010001010100100100000000000",--20823
"111110010000000010010100000000000000",--20824
"001101001000000001100000000000000011",--20825
"011100001101000000000000000000000011",--20826
"101110010001111000000001100000000000",--20827
"011111001011000000110000000000010000",--20828
"000101000000000000000101000101101100",--20829
"111110001000001001010100100000000000",--20830
"001101001000000001100000000000001001",--20831
"001111001100000010100000000000000000",--20832
"111110010010001010100100100000000000",--20833
"111110010000000010010100000000000000",--20834
"111110001010001000110010100000000000",--20835
"001111001100000010010000000000000001",--20836
"111110001010001010010010100000000000",--20837
"111110010000000001010010100000000000",--20838
"111110000110001001000001100000000000",--20839
"001111001100000001000000000000000010",--20840
"111110000110001001000001100000000000",--20841
"111110001010000000110001100000000000",--20842
"011111001011000000110000000000000001",--20843
"111110000110010000010001100000000000",--20844
"111110001110001001110010000000000000",--20845
"111110001100001000110001100000000000",--20846
"111110001000010000110001100000000000",--20847
"010110000111000000000000000000011001",--20848
"001101001000000001000000000000000110",--20849
"011100001001000000000000000000000110",--20850
"111110000110100000000001100000000000",--20851
"111110001110010000110001100000000000",--20852
"001111000110000001000000000000000100",--20853
"111110000110001001000001100000000000",--20854
"001011000000000000110000000100101111",--20855
"000101000000000000000101000101111110",--20856
"111110000110100000000001100000000000",--20857
"111110001110000000110001100000000000",--20858
"001111000110000001000000000000000100",--20859
"111110000110001001000001100000000000",--20860
"001011000000000000110000000100101111",--20861
"001111000000000000110000000100101111",--20862
"101111001001110001001011110111001100",--20863
"101111001001100001001100110011001101",--20864
"010110001001000000110000000000001000",--20865
"101000000011111000000001000000000000",--20866
"101001000000000000010000000000000001",--20867
"001001111100000111111111111111111000",--20868
"101001111100010111100000000000001001",--20869
"000111000000000000000000110101111110",--20870
"101001111100000111100000000000001001",--20871
"001101111100000111111111111111111000",--20872
"011100000011000000000000000000001001",--20873
"101001000000000000010000000000000001",--20874
"001101111100000000101111111111111001",--20875
"001001111100000111111111111111111000",--20876
"101001111100010111100000000000001001",--20877
"000111000000000000000000111111111011",--20878
"101001111100000111100000000000001001",--20879
"001101111100000111111111111111111000",--20880
"011100000011000000000000000000110110",--20881
"000101000000000000000101000110100010",--20882
"101001000000000000010000000000000001",--20883
"001101111100000000101111111111111010",--20884
"001001111100000111111111111111111000",--20885
"101001111100010111100000000000001001",--20886
"000111000000000000000000110101111110",--20887
"101001111100000111100000000000001001",--20888
"001101111100000111111111111111111000",--20889
"011100000011000000000000000000101101",--20890
"101001000000000000010000000000000001",--20891
"001101111100000000101111111111111001",--20892
"101001111100010111100000000000001001",--20893
"000111000000000000000000111111111011",--20894
"101001111100000111100000000000001001",--20895
"001101111100000111111111111111111000",--20896
"011100000011000000000000000000100110",--20897
"101111000111110000110011101111011010",--20898
"101111000111100000110111010000001101",--20899
"001111111100000001001111111111111101",--20900
"111110001000001000110001100000000000",--20901
"001111000000000001000000000100100110",--20902
"001111000000000001010000000101100100",--20903
"111110001000001001010010000000000000",--20904
"001111000000000001010000000100100111",--20905
"001111000000000001100000000101100101",--20906
"111110001010001001100010100000000000",--20907
"111110001000000001010010000000000000",--20908
"001111000000000001010000000100101000",--20909
"001111000000000001100000000101100110",--20910
"111110001010001001100010100000000000",--20911
"111110001000000001010010000000000010",--20912
"010110001001000000000000000000000001",--20913
"000101000000000000000101000110110100",--20914
"101110000001111000000010000000000000",--20915
"111110000110001001000001100000000000",--20916
"001101111100000000011111111111111011",--20917
"001101000010000000010000000000000111",--20918
"001111000010000001000000000000000000",--20919
"111110000110001001000001100000000000",--20920
"001111000000000001000000000100100000",--20921
"001111000000000001010000000100100011",--20922
"111110000110001001010010100000000000",--20923
"111110001000000001010010000000000000",--20924
"001011000000000001000000000100100000",--20925
"001111000000000001000000000100100001",--20926
"001111000000000001010000000100100100",--20927
"111110000110001001010010100000000000",--20928
"111110001000000001010010000000000000",--20929
"001011000000000001000000000100100001",--20930
"001111000000000001000000000100100010",--20931
"001111000000000001010000000100100101",--20932
"111110000110001001010001100000000000",--20933
"111110001000000000110001100000000000",--20934
"001011000000000000110000000100100010",--20935
"101001000000000001000000000001110100",--20936
"001101111100000000011111111111111110",--20937
"001101111100000000101111111111111111",--20938
"001101111100000000110000000000000000",--20939
"000101000000000000000100000011011011",--20940
"001001111100000000100000000000000000",--20941
"001001111100000000111111111111111111",--20942
"001001111100000000011111111111111110",--20943
"010000000011000000000000000011101011",--20944
"001101000000000001000000000011111110",--20945
"001111000110000000110000000000000000",--20946
"001011000000000000110000000100010010",--20947
"001111000110000000110000000000000001",--20948
"001011000000000000110000000100010011",--20949
"001111000110000000110000000000000010",--20950
"001011000000000000110000000100010100",--20951
"001101000000000001010000000110101010",--20952
"101001001010010001010000000000000001",--20953
"001001111100000001001111111111111101",--20954
"010111001011000000000000000011010111",--20955
"001101001010000001100000000101101101",--20956
"001101001100000001110000000000001010",--20957
"001101001100000010000000000000000001",--20958
"001111000110000000110000000000000000",--20959
"001101001100000010010000000000000101",--20960
"001111010010000001000000000000000000",--20961
"111110000110010001000001100000000000",--20962
"001011001110000000110000000000000000",--20963
"001111000110000000110000000000000001",--20964
"001111010010000001000000000000000001",--20965
"111110000110010001000001100000000000",--20966
"001011001110000000110000000000000001",--20967
"001111000110000000110000000000000010",--20968
"001111010010000001000000000000000010",--20969
"111110000110010001000001100000000000",--20970
"001011001110000000110000000000000010",--20971
"011111010001000000100000000000001110",--20972
"001101001100000001100000000000000100",--20973
"001111001110000000110000000000000000",--20974
"001111001110000001000000000000000001",--20975
"001111001110000001010000000000000010",--20976
"001111001100000001100000000000000000",--20977
"111110001100001000110001100000000000",--20978
"001111001100000001100000000000000001",--20979
"111110001100001001000010000000000000",--20980
"111110000110000001000001100000000000",--20981
"001111001100000001000000000000000010",--20982
"111110001000001001010010000000000000",--20983
"111110000110000001000001100000000000",--20984
"001011001110000000110000000000000011",--20985
"000101000000000000000101001000100000",--20986
"010111010001000000100000000000100100",--20987
"001111001110000000110000000000000000",--20988
"001111001110000001000000000000000001",--20989
"001111001110000001010000000000000010",--20990
"111110000110001000110011000000000000",--20991
"001101001100000010010000000000000100",--20992
"001111010010000001110000000000000000",--20993
"111110001100001001110011000000000000",--20994
"111110001000001001000011100000000000",--20995
"001111010010000010000000000000000001",--20996
"111110001110001010000011100000000000",--20997
"111110001100000001110011000000000000",--20998
"111110001010001001010011100000000000",--20999
"001111010010000010000000000000000010",--21000
"111110001110001010000011100000000000",--21001
"111110001100000001110011000000000000",--21002
"001101001100000010010000000000000011",--21003
"011100010011000000000000000000000011",--21004
"101110001101111000000001100000000000",--21005
"011111010001000000110000000000010000",--21006
"000101000000000000000101001000011110",--21007
"111110001000001001010011100000000000",--21008
"001101001100000001100000000000001001",--21009
"001111001100000010000000000000000000",--21010
"111110001110001010000011100000000000",--21011
"111110001100000001110011000000000000",--21012
"111110001010001000110010100000000000",--21013
"001111001100000001110000000000000001",--21014
"111110001010001001110010100000000000",--21015
"111110001100000001010010100000000000",--21016
"111110000110001001000001100000000000",--21017
"001111001100000001000000000000000010",--21018
"111110000110001001000001100000000000",--21019
"111110001010000000110001100000000000",--21020
"011111010001000000110000000000000001",--21021
"111110000110010000010001100000000000",--21022
"001011001110000000110000000000000011",--21023
"101001001010010001010000000000000001",--21024
"010111001011000000000000000010010001",--21025
"001101001010000001100000000101101101",--21026
"001101001100000001110000000000001010",--21027
"001101001100000010000000000000000001",--21028
"001111000110000000110000000000000000",--21029
"001101001100000010010000000000000101",--21030
"001111010010000001000000000000000000",--21031
"111110000110010001000001100000000000",--21032
"001011001110000000110000000000000000",--21033
"001111000110000000110000000000000001",--21034
"001111010010000001000000000000000001",--21035
"111110000110010001000001100000000000",--21036
"001011001110000000110000000000000001",--21037
"001111000110000000110000000000000010",--21038
"001111010010000001000000000000000010",--21039
"111110000110010001000001100000000000",--21040
"001011001110000000110000000000000010",--21041
"011111010001000000100000000000001110",--21042
"001101001100000001100000000000000100",--21043
"001111001110000000110000000000000000",--21044
"001111001110000001000000000000000001",--21045
"001111001110000001010000000000000010",--21046
"001111001100000001100000000000000000",--21047
"111110001100001000110001100000000000",--21048
"001111001100000001100000000000000001",--21049
"111110001100001001000010000000000000",--21050
"111110000110000001000001100000000000",--21051
"001111001100000001000000000000000010",--21052
"111110001000001001010010000000000000",--21053
"111110000110000001000001100000000000",--21054
"001011001110000000110000000000000011",--21055
"000101000000000000000101001001100110",--21056
"010111010001000000100000000000100100",--21057
"001111001110000000110000000000000000",--21058
"001111001110000001000000000000000001",--21059
"001111001110000001010000000000000010",--21060
"111110000110001000110011000000000000",--21061
"001101001100000010010000000000000100",--21062
"001111010010000001110000000000000000",--21063
"111110001100001001110011000000000000",--21064
"111110001000001001000011100000000000",--21065
"001111010010000010000000000000000001",--21066
"111110001110001010000011100000000000",--21067
"111110001100000001110011000000000000",--21068
"111110001010001001010011100000000000",--21069
"001111010010000010000000000000000010",--21070
"111110001110001010000011100000000000",--21071
"111110001100000001110011000000000000",--21072
"001101001100000010010000000000000011",--21073
"011100010011000000000000000000000011",--21074
"101110001101111000000001100000000000",--21075
"011111010001000000110000000000010000",--21076
"000101000000000000000101001001100100",--21077
"111110001000001001010011100000000000",--21078
"001101001100000001100000000000001001",--21079
"001111001100000010000000000000000000",--21080
"111110001110001010000011100000000000",--21081
"111110001100000001110011000000000000",--21082
"111110001010001000110010100000000000",--21083
"001111001100000001110000000000000001",--21084
"111110001010001001110010100000000000",--21085
"111110001100000001010010100000000000",--21086
"111110000110001001000001100000000000",--21087
"001111001100000001000000000000000010",--21088
"111110000110001001000001100000000000",--21089
"111110001010000000110001100000000000",--21090
"011111010001000000110000000000000001",--21091
"111110000110010000010001100000000000",--21092
"001011001110000000110000000000000011",--21093
"101001001010010001010000000000000001",--21094
"010111001011000000000000000001001011",--21095
"001101001010000001100000000101101101",--21096
"001101001100000001110000000000001010",--21097
"001101001100000010000000000000000001",--21098
"001111000110000000110000000000000000",--21099
"001101001100000010010000000000000101",--21100
"001111010010000001000000000000000000",--21101
"111110000110010001000001100000000000",--21102
"001011001110000000110000000000000000",--21103
"001111000110000000110000000000000001",--21104
"001111010010000001000000000000000001",--21105
"111110000110010001000001100000000000",--21106
"001011001110000000110000000000000001",--21107
"001111000110000000110000000000000010",--21108
"001111010010000001000000000000000010",--21109
"111110000110010001000001100000000000",--21110
"001011001110000000110000000000000010",--21111
"011111010001000000100000000000001110",--21112
"001101001100000001100000000000000100",--21113
"001111001110000000110000000000000000",--21114
"001111001110000001000000000000000001",--21115
"001111001110000001010000000000000010",--21116
"001111001100000001100000000000000000",--21117
"111110001100001000110001100000000000",--21118
"001111001100000001100000000000000001",--21119
"111110001100001001000010000000000000",--21120
"111110000110000001000001100000000000",--21121
"001111001100000001000000000000000010",--21122
"111110001000001001010010000000000000",--21123
"111110000110000001000001100000000000",--21124
"001011001110000000110000000000000011",--21125
"000101000000000000000101001010101100",--21126
"010111010001000000100000000000100100",--21127
"001111001110000000110000000000000000",--21128
"001111001110000001000000000000000001",--21129
"001111001110000001010000000000000010",--21130
"111110000110001000110011000000000000",--21131
"001101001100000010010000000000000100",--21132
"001111010010000001110000000000000000",--21133
"111110001100001001110011000000000000",--21134
"111110001000001001000011100000000000",--21135
"001111010010000010000000000000000001",--21136
"111110001110001010000011100000000000",--21137
"111110001100000001110011000000000000",--21138
"111110001010001001010011100000000000",--21139
"001111010010000010000000000000000010",--21140
"111110001110001010000011100000000000",--21141
"111110001100000001110011000000000000",--21142
"001101001100000010010000000000000011",--21143
"011100010011000000000000000000000011",--21144
"101110001101111000000001100000000000",--21145
"011111010001000000110000000000010000",--21146
"000101000000000000000101001010101010",--21147
"111110001000001001010011100000000000",--21148
"001101001100000001100000000000001001",--21149
"001111001100000010000000000000000000",--21150
"111110001110001010000011100000000000",--21151
"111110001100000001110011000000000000",--21152
"111110001010001000110010100000000000",--21153
"001111001100000001110000000000000001",--21154
"111110001010001001110010100000000000",--21155
"111110001100000001010010100000000000",--21156
"111110000110001001000001100000000000",--21157
"001111001100000001000000000000000010",--21158
"111110000110001001000001100000000000",--21159
"111110001010000000110001100000000000",--21160
"011111010001000000110000000000000001",--21161
"111110000110010000010001100000000000",--21162
"001011001110000000110000000000000011",--21163
"101001001010010000100000000000000001",--21164
"101000000111111000000000100000000000",--21165
"001001111100000111111111111111111100",--21166
"101001111100010111100000000000000101",--21167
"000111000000000000000000011001101110",--21168
"101001111100000111100000000000000101",--21169
"001101111100000111111111111111111100",--21170
"101001000000000001000000000001110110",--21171
"001101111100000000011111111111111101",--21172
"001101111100000000100000000000000000",--21173
"001101111100000000111111111111111111",--21174
"001001111100000111111111111111111100",--21175
"101001111100010111100000000000000101",--21176
"000111000000000000000100000011011010",--21177
"101001111100000111100000000000000101",--21178
"001101111100000111111111111111111100",--21179
"001101111100000000011111111111111110",--21180
"010011000011000000010000000011101100",--21181
"001101000000000000100000000011111111",--21182
"001101111100000000111111111111111111",--21183
"001111000110000000110000000000000000",--21184
"001011000000000000110000000100010010",--21185
"001111000110000000110000000000000001",--21186
"001011000000000000110000000100010011",--21187
"001111000110000000110000000000000010",--21188
"001011000000000000110000000100010100",--21189
"001101000000000001000000000110101010",--21190
"101001001000010001000000000000000001",--21191
"001001111100000000101111111111111101",--21192
"010111001001000000000000000011010111",--21193
"001101001000000001010000000101101101",--21194
"001101001010000001100000000000001010",--21195
"001101001010000001110000000000000001",--21196
"001111000110000000110000000000000000",--21197
"001101001010000010000000000000000101",--21198
"001111010000000001000000000000000000",--21199
"111110000110010001000001100000000000",--21200
"001011001100000000110000000000000000",--21201
"001111000110000000110000000000000001",--21202
"001111010000000001000000000000000001",--21203
"111110000110010001000001100000000000",--21204
"001011001100000000110000000000000001",--21205
"001111000110000000110000000000000010",--21206
"001111010000000001000000000000000010",--21207
"111110000110010001000001100000000000",--21208
"001011001100000000110000000000000010",--21209
"011111001111000000100000000000001110",--21210
"001101001010000001010000000000000100",--21211
"001111001100000000110000000000000000",--21212
"001111001100000001000000000000000001",--21213
"001111001100000001010000000000000010",--21214
"001111001010000001100000000000000000",--21215
"111110001100001000110001100000000000",--21216
"001111001010000001100000000000000001",--21217
"111110001100001001000010000000000000",--21218
"111110000110000001000001100000000000",--21219
"001111001010000001000000000000000010",--21220
"111110001000001001010010000000000000",--21221
"111110000110000001000001100000000000",--21222
"001011001100000000110000000000000011",--21223
"000101000000000000000101001100001110",--21224
"010111001111000000100000000000100100",--21225
"001111001100000000110000000000000000",--21226
"001111001100000001000000000000000001",--21227
"001111001100000001010000000000000010",--21228
"111110000110001000110011000000000000",--21229
"001101001010000010000000000000000100",--21230
"001111010000000001110000000000000000",--21231
"111110001100001001110011000000000000",--21232
"111110001000001001000011100000000000",--21233
"001111010000000010000000000000000001",--21234
"111110001110001010000011100000000000",--21235
"111110001100000001110011000000000000",--21236
"111110001010001001010011100000000000",--21237
"001111010000000010000000000000000010",--21238
"111110001110001010000011100000000000",--21239
"111110001100000001110011000000000000",--21240
"001101001010000010000000000000000011",--21241
"011100010001000000000000000000000011",--21242
"101110001101111000000001100000000000",--21243
"011111001111000000110000000000010000",--21244
"000101000000000000000101001100001100",--21245
"111110001000001001010011100000000000",--21246
"001101001010000001010000000000001001",--21247
"001111001010000010000000000000000000",--21248
"111110001110001010000011100000000000",--21249
"111110001100000001110011000000000000",--21250
"111110001010001000110010100000000000",--21251
"001111001010000001110000000000000001",--21252
"111110001010001001110010100000000000",--21253
"111110001100000001010010100000000000",--21254
"111110000110001001000001100000000000",--21255
"001111001010000001000000000000000010",--21256
"111110000110001001000001100000000000",--21257
"111110001010000000110001100000000000",--21258
"011111001111000000110000000000000001",--21259
"111110000110010000010001100000000000",--21260
"001011001100000000110000000000000011",--21261
"101001001000010001000000000000000001",--21262
"010111001001000000000000000010010001",--21263
"001101001000000001010000000101101101",--21264
"001101001010000001100000000000001010",--21265
"001101001010000001110000000000000001",--21266
"001111000110000000110000000000000000",--21267
"001101001010000010000000000000000101",--21268
"001111010000000001000000000000000000",--21269
"111110000110010001000001100000000000",--21270
"001011001100000000110000000000000000",--21271
"001111000110000000110000000000000001",--21272
"001111010000000001000000000000000001",--21273
"111110000110010001000001100000000000",--21274
"001011001100000000110000000000000001",--21275
"001111000110000000110000000000000010",--21276
"001111010000000001000000000000000010",--21277
"111110000110010001000001100000000000",--21278
"001011001100000000110000000000000010",--21279
"011111001111000000100000000000001110",--21280
"001101001010000001010000000000000100",--21281
"001111001100000000110000000000000000",--21282
"001111001100000001000000000000000001",--21283
"001111001100000001010000000000000010",--21284
"001111001010000001100000000000000000",--21285
"111110001100001000110001100000000000",--21286
"001111001010000001100000000000000001",--21287
"111110001100001001000010000000000000",--21288
"111110000110000001000001100000000000",--21289
"001111001010000001000000000000000010",--21290
"111110001000001001010010000000000000",--21291
"111110000110000001000001100000000000",--21292
"001011001100000000110000000000000011",--21293
"000101000000000000000101001101010100",--21294
"010111001111000000100000000000100100",--21295
"001111001100000000110000000000000000",--21296
"001111001100000001000000000000000001",--21297
"001111001100000001010000000000000010",--21298
"111110000110001000110011000000000000",--21299
"001101001010000010000000000000000100",--21300
"001111010000000001110000000000000000",--21301
"111110001100001001110011000000000000",--21302
"111110001000001001000011100000000000",--21303
"001111010000000010000000000000000001",--21304
"111110001110001010000011100000000000",--21305
"111110001100000001110011000000000000",--21306
"111110001010001001010011100000000000",--21307
"001111010000000010000000000000000010",--21308
"111110001110001010000011100000000000",--21309
"111110001100000001110011000000000000",--21310
"001101001010000010000000000000000011",--21311
"011100010001000000000000000000000011",--21312
"101110001101111000000001100000000000",--21313
"011111001111000000110000000000010000",--21314
"000101000000000000000101001101010010",--21315
"111110001000001001010011100000000000",--21316
"001101001010000001010000000000001001",--21317
"001111001010000010000000000000000000",--21318
"111110001110001010000011100000000000",--21319
"111110001100000001110011000000000000",--21320
"111110001010001000110010100000000000",--21321
"001111001010000001110000000000000001",--21322
"111110001010001001110010100000000000",--21323
"111110001100000001010010100000000000",--21324
"111110000110001001000001100000000000",--21325
"001111001010000001000000000000000010",--21326
"111110000110001001000001100000000000",--21327
"111110001010000000110001100000000000",--21328
"011111001111000000110000000000000001",--21329
"111110000110010000010001100000000000",--21330
"001011001100000000110000000000000011",--21331
"101001001000010001000000000000000001",--21332
"010111001001000000000000000001001011",--21333
"001101001000000001010000000101101101",--21334
"001101001010000001100000000000001010",--21335
"001101001010000001110000000000000001",--21336
"001111000110000000110000000000000000",--21337
"001101001010000010000000000000000101",--21338
"001111010000000001000000000000000000",--21339
"111110000110010001000001100000000000",--21340
"001011001100000000110000000000000000",--21341
"001111000110000000110000000000000001",--21342
"001111010000000001000000000000000001",--21343
"111110000110010001000001100000000000",--21344
"001011001100000000110000000000000001",--21345
"001111000110000000110000000000000010",--21346
"001111010000000001000000000000000010",--21347
"111110000110010001000001100000000000",--21348
"001011001100000000110000000000000010",--21349
"011111001111000000100000000000001110",--21350
"001101001010000001010000000000000100",--21351
"001111001100000000110000000000000000",--21352
"001111001100000001000000000000000001",--21353
"001111001100000001010000000000000010",--21354
"001111001010000001100000000000000000",--21355
"111110001100001000110001100000000000",--21356
"001111001010000001100000000000000001",--21357
"111110001100001001000010000000000000",--21358
"111110000110000001000001100000000000",--21359
"001111001010000001000000000000000010",--21360
"111110001000001001010010000000000000",--21361
"111110000110000001000001100000000000",--21362
"001011001100000000110000000000000011",--21363
"000101000000000000000101001110011010",--21364
"010111001111000000100000000000100100",--21365
"001111001100000000110000000000000000",--21366
"001111001100000001000000000000000001",--21367
"001111001100000001010000000000000010",--21368
"111110000110001000110011000000000000",--21369
"001101001010000010000000000000000100",--21370
"001111010000000001110000000000000000",--21371
"111110001100001001110011000000000000",--21372
"111110001000001001000011100000000000",--21373
"001111010000000010000000000000000001",--21374
"111110001110001010000011100000000000",--21375
"111110001100000001110011000000000000",--21376
"111110001010001001010011100000000000",--21377
"001111010000000010000000000000000010",--21378
"111110001110001010000011100000000000",--21379
"111110001100000001110011000000000000",--21380
"001101001010000010000000000000000011",--21381
"011100010001000000000000000000000011",--21382
"101110001101111000000001100000000000",--21383
"011111001111000000110000000000010000",--21384
"000101000000000000000101001110011000",--21385
"111110001000001001010011100000000000",--21386
"001101001010000001010000000000001001",--21387
"001111001010000010000000000000000000",--21388
"111110001110001010000011100000000000",--21389
"111110001100000001110011000000000000",--21390
"111110001010001000110010100000000000",--21391
"001111001010000001110000000000000001",--21392
"111110001010001001110010100000000000",--21393
"111110001100000001010010100000000000",--21394
"111110000110001001000001100000000000",--21395
"001111001010000001000000000000000010",--21396
"111110000110001001000001100000000000",--21397
"111110001010000000110001100000000000",--21398
"011111001111000000110000000000000001",--21399
"111110000110010000010001100000000000",--21400
"001011001100000000110000000000000011",--21401
"101001001000010000100000000000000001",--21402
"101000000111111000000000100000000000",--21403
"001001111100000111111111111111111100",--21404
"101001111100010111100000000000000101",--21405
"000111000000000000000000011001101110",--21406
"101001111100000111100000000000000101",--21407
"001101111100000111111111111111111100",--21408
"101001000000000001000000000001110110",--21409
"001101111100000000011111111111111101",--21410
"001101111100000000100000000000000000",--21411
"001101111100000000111111111111111111",--21412
"001001111100000111111111111111111100",--21413
"101001111100010111100000000000000101",--21414
"000111000000000000000100000011011010",--21415
"101001111100000111100000000000000101",--21416
"001101111100000111111111111111111100",--21417
"001101111100000000011111111111111110",--21418
"010011000011000000100000000011101100",--21419
"001101000000000000100000000100000000",--21420
"001101111100000000111111111111111111",--21421
"001111000110000000110000000000000000",--21422
"001011000000000000110000000100010010",--21423
"001111000110000000110000000000000001",--21424
"001011000000000000110000000100010011",--21425
"001111000110000000110000000000000010",--21426
"001011000000000000110000000100010100",--21427
"001101000000000001000000000110101010",--21428
"101001001000010001000000000000000001",--21429
"001001111100000000101111111111111101",--21430
"010111001001000000000000000011010111",--21431
"001101001000000001010000000101101101",--21432
"001101001010000001100000000000001010",--21433
"001101001010000001110000000000000001",--21434
"001111000110000000110000000000000000",--21435
"001101001010000010000000000000000101",--21436
"001111010000000001000000000000000000",--21437
"111110000110010001000001100000000000",--21438
"001011001100000000110000000000000000",--21439
"001111000110000000110000000000000001",--21440
"001111010000000001000000000000000001",--21441
"111110000110010001000001100000000000",--21442
"001011001100000000110000000000000001",--21443
"001111000110000000110000000000000010",--21444
"001111010000000001000000000000000010",--21445
"111110000110010001000001100000000000",--21446
"001011001100000000110000000000000010",--21447
"011111001111000000100000000000001110",--21448
"001101001010000001010000000000000100",--21449
"001111001100000000110000000000000000",--21450
"001111001100000001000000000000000001",--21451
"001111001100000001010000000000000010",--21452
"001111001010000001100000000000000000",--21453
"111110001100001000110001100000000000",--21454
"001111001010000001100000000000000001",--21455
"111110001100001001000010000000000000",--21456
"111110000110000001000001100000000000",--21457
"001111001010000001000000000000000010",--21458
"111110001000001001010010000000000000",--21459
"111110000110000001000001100000000000",--21460
"001011001100000000110000000000000011",--21461
"000101000000000000000101001111111100",--21462
"010111001111000000100000000000100100",--21463
"001111001100000000110000000000000000",--21464
"001111001100000001000000000000000001",--21465
"001111001100000001010000000000000010",--21466
"111110000110001000110011000000000000",--21467
"001101001010000010000000000000000100",--21468
"001111010000000001110000000000000000",--21469
"111110001100001001110011000000000000",--21470
"111110001000001001000011100000000000",--21471
"001111010000000010000000000000000001",--21472
"111110001110001010000011100000000000",--21473
"111110001100000001110011000000000000",--21474
"111110001010001001010011100000000000",--21475
"001111010000000010000000000000000010",--21476
"111110001110001010000011100000000000",--21477
"111110001100000001110011000000000000",--21478
"001101001010000010000000000000000011",--21479
"011100010001000000000000000000000011",--21480
"101110001101111000000001100000000000",--21481
"011111001111000000110000000000010000",--21482
"000101000000000000000101001111111010",--21483
"111110001000001001010011100000000000",--21484
"001101001010000001010000000000001001",--21485
"001111001010000010000000000000000000",--21486
"111110001110001010000011100000000000",--21487
"111110001100000001110011000000000000",--21488
"111110001010001000110010100000000000",--21489
"001111001010000001110000000000000001",--21490
"111110001010001001110010100000000000",--21491
"111110001100000001010010100000000000",--21492
"111110000110001001000001100000000000",--21493
"001111001010000001000000000000000010",--21494
"111110000110001001000001100000000000",--21495
"111110001010000000110001100000000000",--21496
"011111001111000000110000000000000001",--21497
"111110000110010000010001100000000000",--21498
"001011001100000000110000000000000011",--21499
"101001001000010001000000000000000001",--21500
"010111001001000000000000000010010001",--21501
"001101001000000001010000000101101101",--21502
"001101001010000001100000000000001010",--21503
"001101001010000001110000000000000001",--21504
"001111000110000000110000000000000000",--21505
"001101001010000010000000000000000101",--21506
"001111010000000001000000000000000000",--21507
"111110000110010001000001100000000000",--21508
"001011001100000000110000000000000000",--21509
"001111000110000000110000000000000001",--21510
"001111010000000001000000000000000001",--21511
"111110000110010001000001100000000000",--21512
"001011001100000000110000000000000001",--21513
"001111000110000000110000000000000010",--21514
"001111010000000001000000000000000010",--21515
"111110000110010001000001100000000000",--21516
"001011001100000000110000000000000010",--21517
"011111001111000000100000000000001110",--21518
"001101001010000001010000000000000100",--21519
"001111001100000000110000000000000000",--21520
"001111001100000001000000000000000001",--21521
"001111001100000001010000000000000010",--21522
"001111001010000001100000000000000000",--21523
"111110001100001000110001100000000000",--21524
"001111001010000001100000000000000001",--21525
"111110001100001001000010000000000000",--21526
"111110000110000001000001100000000000",--21527
"001111001010000001000000000000000010",--21528
"111110001000001001010010000000000000",--21529
"111110000110000001000001100000000000",--21530
"001011001100000000110000000000000011",--21531
"000101000000000000000101010001000010",--21532
"010111001111000000100000000000100100",--21533
"001111001100000000110000000000000000",--21534
"001111001100000001000000000000000001",--21535
"001111001100000001010000000000000010",--21536
"111110000110001000110011000000000000",--21537
"001101001010000010000000000000000100",--21538
"001111010000000001110000000000000000",--21539
"111110001100001001110011000000000000",--21540
"111110001000001001000011100000000000",--21541
"001111010000000010000000000000000001",--21542
"111110001110001010000011100000000000",--21543
"111110001100000001110011000000000000",--21544
"111110001010001001010011100000000000",--21545
"001111010000000010000000000000000010",--21546
"111110001110001010000011100000000000",--21547
"111110001100000001110011000000000000",--21548
"001101001010000010000000000000000011",--21549
"011100010001000000000000000000000011",--21550
"101110001101111000000001100000000000",--21551
"011111001111000000110000000000010000",--21552
"000101000000000000000101010001000000",--21553
"111110001000001001010011100000000000",--21554
"001101001010000001010000000000001001",--21555
"001111001010000010000000000000000000",--21556
"111110001110001010000011100000000000",--21557
"111110001100000001110011000000000000",--21558
"111110001010001000110010100000000000",--21559
"001111001010000001110000000000000001",--21560
"111110001010001001110010100000000000",--21561
"111110001100000001010010100000000000",--21562
"111110000110001001000001100000000000",--21563
"001111001010000001000000000000000010",--21564
"111110000110001001000001100000000000",--21565
"111110001010000000110001100000000000",--21566
"011111001111000000110000000000000001",--21567
"111110000110010000010001100000000000",--21568
"001011001100000000110000000000000011",--21569
"101001001000010001000000000000000001",--21570
"010111001001000000000000000001001011",--21571
"001101001000000001010000000101101101",--21572
"001101001010000001100000000000001010",--21573
"001101001010000001110000000000000001",--21574
"001111000110000000110000000000000000",--21575
"001101001010000010000000000000000101",--21576
"001111010000000001000000000000000000",--21577
"111110000110010001000001100000000000",--21578
"001011001100000000110000000000000000",--21579
"001111000110000000110000000000000001",--21580
"001111010000000001000000000000000001",--21581
"111110000110010001000001100000000000",--21582
"001011001100000000110000000000000001",--21583
"001111000110000000110000000000000010",--21584
"001111010000000001000000000000000010",--21585
"111110000110010001000001100000000000",--21586
"001011001100000000110000000000000010",--21587
"011111001111000000100000000000001110",--21588
"001101001010000001010000000000000100",--21589
"001111001100000000110000000000000000",--21590
"001111001100000001000000000000000001",--21591
"001111001100000001010000000000000010",--21592
"001111001010000001100000000000000000",--21593
"111110001100001000110001100000000000",--21594
"001111001010000001100000000000000001",--21595
"111110001100001001000010000000000000",--21596
"111110000110000001000001100000000000",--21597
"001111001010000001000000000000000010",--21598
"111110001000001001010010000000000000",--21599
"111110000110000001000001100000000000",--21600
"001011001100000000110000000000000011",--21601
"000101000000000000000101010010001000",--21602
"010111001111000000100000000000100100",--21603
"001111001100000000110000000000000000",--21604
"001111001100000001000000000000000001",--21605
"001111001100000001010000000000000010",--21606
"111110000110001000110011000000000000",--21607
"001101001010000010000000000000000100",--21608
"001111010000000001110000000000000000",--21609
"111110001100001001110011000000000000",--21610
"111110001000001001000011100000000000",--21611
"001111010000000010000000000000000001",--21612
"111110001110001010000011100000000000",--21613
"111110001100000001110011000000000000",--21614
"111110001010001001010011100000000000",--21615
"001111010000000010000000000000000010",--21616
"111110001110001010000011100000000000",--21617
"111110001100000001110011000000000000",--21618
"001101001010000010000000000000000011",--21619
"011100010001000000000000000000000011",--21620
"101110001101111000000001100000000000",--21621
"011111001111000000110000000000010000",--21622
"000101000000000000000101010010000110",--21623
"111110001000001001010011100000000000",--21624
"001101001010000001010000000000001001",--21625
"001111001010000010000000000000000000",--21626
"111110001110001010000011100000000000",--21627
"111110001100000001110011000000000000",--21628
"111110001010001000110010100000000000",--21629
"001111001010000001110000000000000001",--21630
"111110001010001001110010100000000000",--21631
"111110001100000001010010100000000000",--21632
"111110000110001001000001100000000000",--21633
"001111001010000001000000000000000010",--21634
"111110000110001001000001100000000000",--21635
"111110001010000000110001100000000000",--21636
"011111001111000000110000000000000001",--21637
"111110000110010000010001100000000000",--21638
"001011001100000000110000000000000011",--21639
"101001001000010000100000000000000001",--21640
"101000000111111000000000100000000000",--21641
"001001111100000111111111111111111100",--21642
"101001111100010111100000000000000101",--21643
"000111000000000000000000011001101110",--21644
"101001111100000111100000000000000101",--21645
"001101111100000111111111111111111100",--21646
"101001000000000001000000000001110110",--21647
"001101111100000000011111111111111101",--21648
"001101111100000000100000000000000000",--21649
"001101111100000000111111111111111111",--21650
"001001111100000111111111111111111100",--21651
"101001111100010111100000000000000101",--21652
"000111000000000000000100000011011010",--21653
"101001111100000111100000000000000101",--21654
"001101111100000111111111111111111100",--21655
"001101111100000000011111111111111110",--21656
"010011000011000000110000000011101100",--21657
"001101000000000000100000000100000001",--21658
"001101111100000000111111111111111111",--21659
"001111000110000000110000000000000000",--21660
"001011000000000000110000000100010010",--21661
"001111000110000000110000000000000001",--21662
"001011000000000000110000000100010011",--21663
"001111000110000000110000000000000010",--21664
"001011000000000000110000000100010100",--21665
"001101000000000001000000000110101010",--21666
"101001001000010001000000000000000001",--21667
"001001111100000000101111111111111101",--21668
"010111001001000000000000000011010111",--21669
"001101001000000001010000000101101101",--21670
"001101001010000001100000000000001010",--21671
"001101001010000001110000000000000001",--21672
"001111000110000000110000000000000000",--21673
"001101001010000010000000000000000101",--21674
"001111010000000001000000000000000000",--21675
"111110000110010001000001100000000000",--21676
"001011001100000000110000000000000000",--21677
"001111000110000000110000000000000001",--21678
"001111010000000001000000000000000001",--21679
"111110000110010001000001100000000000",--21680
"001011001100000000110000000000000001",--21681
"001111000110000000110000000000000010",--21682
"001111010000000001000000000000000010",--21683
"111110000110010001000001100000000000",--21684
"001011001100000000110000000000000010",--21685
"011111001111000000100000000000001110",--21686
"001101001010000001010000000000000100",--21687
"001111001100000000110000000000000000",--21688
"001111001100000001000000000000000001",--21689
"001111001100000001010000000000000010",--21690
"001111001010000001100000000000000000",--21691
"111110001100001000110001100000000000",--21692
"001111001010000001100000000000000001",--21693
"111110001100001001000010000000000000",--21694
"111110000110000001000001100000000000",--21695
"001111001010000001000000000000000010",--21696
"111110001000001001010010000000000000",--21697
"111110000110000001000001100000000000",--21698
"001011001100000000110000000000000011",--21699
"000101000000000000000101010011101010",--21700
"010111001111000000100000000000100100",--21701
"001111001100000000110000000000000000",--21702
"001111001100000001000000000000000001",--21703
"001111001100000001010000000000000010",--21704
"111110000110001000110011000000000000",--21705
"001101001010000010000000000000000100",--21706
"001111010000000001110000000000000000",--21707
"111110001100001001110011000000000000",--21708
"111110001000001001000011100000000000",--21709
"001111010000000010000000000000000001",--21710
"111110001110001010000011100000000000",--21711
"111110001100000001110011000000000000",--21712
"111110001010001001010011100000000000",--21713
"001111010000000010000000000000000010",--21714
"111110001110001010000011100000000000",--21715
"111110001100000001110011000000000000",--21716
"001101001010000010000000000000000011",--21717
"011100010001000000000000000000000011",--21718
"101110001101111000000001100000000000",--21719
"011111001111000000110000000000010000",--21720
"000101000000000000000101010011101000",--21721
"111110001000001001010011100000000000",--21722
"001101001010000001010000000000001001",--21723
"001111001010000010000000000000000000",--21724
"111110001110001010000011100000000000",--21725
"111110001100000001110011000000000000",--21726
"111110001010001000110010100000000000",--21727
"001111001010000001110000000000000001",--21728
"111110001010001001110010100000000000",--21729
"111110001100000001010010100000000000",--21730
"111110000110001001000001100000000000",--21731
"001111001010000001000000000000000010",--21732
"111110000110001001000001100000000000",--21733
"111110001010000000110001100000000000",--21734
"011111001111000000110000000000000001",--21735
"111110000110010000010001100000000000",--21736
"001011001100000000110000000000000011",--21737
"101001001000010001000000000000000001",--21738
"010111001001000000000000000010010001",--21739
"001101001000000001010000000101101101",--21740
"001101001010000001100000000000001010",--21741
"001101001010000001110000000000000001",--21742
"001111000110000000110000000000000000",--21743
"001101001010000010000000000000000101",--21744
"001111010000000001000000000000000000",--21745
"111110000110010001000001100000000000",--21746
"001011001100000000110000000000000000",--21747
"001111000110000000110000000000000001",--21748
"001111010000000001000000000000000001",--21749
"111110000110010001000001100000000000",--21750
"001011001100000000110000000000000001",--21751
"001111000110000000110000000000000010",--21752
"001111010000000001000000000000000010",--21753
"111110000110010001000001100000000000",--21754
"001011001100000000110000000000000010",--21755
"011111001111000000100000000000001110",--21756
"001101001010000001010000000000000100",--21757
"001111001100000000110000000000000000",--21758
"001111001100000001000000000000000001",--21759
"001111001100000001010000000000000010",--21760
"001111001010000001100000000000000000",--21761
"111110001100001000110001100000000000",--21762
"001111001010000001100000000000000001",--21763
"111110001100001001000010000000000000",--21764
"111110000110000001000001100000000000",--21765
"001111001010000001000000000000000010",--21766
"111110001000001001010010000000000000",--21767
"111110000110000001000001100000000000",--21768
"001011001100000000110000000000000011",--21769
"000101000000000000000101010100110000",--21770
"010111001111000000100000000000100100",--21771
"001111001100000000110000000000000000",--21772
"001111001100000001000000000000000001",--21773
"001111001100000001010000000000000010",--21774
"111110000110001000110011000000000000",--21775
"001101001010000010000000000000000100",--21776
"001111010000000001110000000000000000",--21777
"111110001100001001110011000000000000",--21778
"111110001000001001000011100000000000",--21779
"001111010000000010000000000000000001",--21780
"111110001110001010000011100000000000",--21781
"111110001100000001110011000000000000",--21782
"111110001010001001010011100000000000",--21783
"001111010000000010000000000000000010",--21784
"111110001110001010000011100000000000",--21785
"111110001100000001110011000000000000",--21786
"001101001010000010000000000000000011",--21787
"011100010001000000000000000000000011",--21788
"101110001101111000000001100000000000",--21789
"011111001111000000110000000000010000",--21790
"000101000000000000000101010100101110",--21791
"111110001000001001010011100000000000",--21792
"001101001010000001010000000000001001",--21793
"001111001010000010000000000000000000",--21794
"111110001110001010000011100000000000",--21795
"111110001100000001110011000000000000",--21796
"111110001010001000110010100000000000",--21797
"001111001010000001110000000000000001",--21798
"111110001010001001110010100000000000",--21799
"111110001100000001010010100000000000",--21800
"111110000110001001000001100000000000",--21801
"001111001010000001000000000000000010",--21802
"111110000110001001000001100000000000",--21803
"111110001010000000110001100000000000",--21804
"011111001111000000110000000000000001",--21805
"111110000110010000010001100000000000",--21806
"001011001100000000110000000000000011",--21807
"101001001000010001000000000000000001",--21808
"010111001001000000000000000001001011",--21809
"001101001000000001010000000101101101",--21810
"001101001010000001100000000000001010",--21811
"001101001010000001110000000000000001",--21812
"001111000110000000110000000000000000",--21813
"001101001010000010000000000000000101",--21814
"001111010000000001000000000000000000",--21815
"111110000110010001000001100000000000",--21816
"001011001100000000110000000000000000",--21817
"001111000110000000110000000000000001",--21818
"001111010000000001000000000000000001",--21819
"111110000110010001000001100000000000",--21820
"001011001100000000110000000000000001",--21821
"001111000110000000110000000000000010",--21822
"001111010000000001000000000000000010",--21823
"111110000110010001000001100000000000",--21824
"001011001100000000110000000000000010",--21825
"011111001111000000100000000000001110",--21826
"001101001010000001010000000000000100",--21827
"001111001100000000110000000000000000",--21828
"001111001100000001000000000000000001",--21829
"001111001100000001010000000000000010",--21830
"001111001010000001100000000000000000",--21831
"111110001100001000110001100000000000",--21832
"001111001010000001100000000000000001",--21833
"111110001100001001000010000000000000",--21834
"111110000110000001000001100000000000",--21835
"001111001010000001000000000000000010",--21836
"111110001000001001010010000000000000",--21837
"111110000110000001000001100000000000",--21838
"001011001100000000110000000000000011",--21839
"000101000000000000000101010101110110",--21840
"010111001111000000100000000000100100",--21841
"001111001100000000110000000000000000",--21842
"001111001100000001000000000000000001",--21843
"001111001100000001010000000000000010",--21844
"111110000110001000110011000000000000",--21845
"001101001010000010000000000000000100",--21846
"001111010000000001110000000000000000",--21847
"111110001100001001110011000000000000",--21848
"111110001000001001000011100000000000",--21849
"001111010000000010000000000000000001",--21850
"111110001110001010000011100000000000",--21851
"111110001100000001110011000000000000",--21852
"111110001010001001010011100000000000",--21853
"001111010000000010000000000000000010",--21854
"111110001110001010000011100000000000",--21855
"111110001100000001110011000000000000",--21856
"001101001010000010000000000000000011",--21857
"011100010001000000000000000000000011",--21858
"101110001101111000000001100000000000",--21859
"011111001111000000110000000000010000",--21860
"000101000000000000000101010101110100",--21861
"111110001000001001010011100000000000",--21862
"001101001010000001010000000000001001",--21863
"001111001010000010000000000000000000",--21864
"111110001110001010000011100000000000",--21865
"111110001100000001110011000000000000",--21866
"111110001010001000110010100000000000",--21867
"001111001010000001110000000000000001",--21868
"111110001010001001110010100000000000",--21869
"111110001100000001010010100000000000",--21870
"111110000110001001000001100000000000",--21871
"001111001010000001000000000000000010",--21872
"111110000110001001000001100000000000",--21873
"111110001010000000110001100000000000",--21874
"011111001111000000110000000000000001",--21875
"111110000110010000010001100000000000",--21876
"001011001100000000110000000000000011",--21877
"101001001000010000100000000000000001",--21878
"101000000111111000000000100000000000",--21879
"001001111100000111111111111111111100",--21880
"101001111100010111100000000000000101",--21881
"000111000000000000000000011001101110",--21882
"101001111100000111100000000000000101",--21883
"001101111100000111111111111111111100",--21884
"101001000000000001000000000001110110",--21885
"001101111100000000011111111111111101",--21886
"001101111100000000100000000000000000",--21887
"001101111100000000111111111111111111",--21888
"001001111100000111111111111111111100",--21889
"101001111100010111100000000000000101",--21890
"000111000000000000000100000011011010",--21891
"101001111100000111100000000000000101",--21892
"001101111100000111111111111111111100",--21893
"001101111100000000011111111111111110",--21894
"010011000010000001001111100000000000",--21895
"001101000000000000010000000100000010",--21896
"001101111100000000111111111111111111",--21897
"001111000110000000110000000000000000",--21898
"001011000000000000110000000100010010",--21899
"001111000110000000110000000000000001",--21900
"001011000000000000110000000100010011",--21901
"001111000110000000110000000000000010",--21902
"001011000000000000110000000100010100",--21903
"001101000000000000100000000110101010",--21904
"101001000100010000100000000000000001",--21905
"001001111100000000011111111111111101",--21906
"010111000101000000000000000011010111",--21907
"001101000100000001000000000101101101",--21908
"001101001000000001010000000000001010",--21909
"001101001000000001100000000000000001",--21910
"001111000110000000110000000000000000",--21911
"001101001000000001110000000000000101",--21912
"001111001110000001000000000000000000",--21913
"111110000110010001000001100000000000",--21914
"001011001010000000110000000000000000",--21915
"001111000110000000110000000000000001",--21916
"001111001110000001000000000000000001",--21917
"111110000110010001000001100000000000",--21918
"001011001010000000110000000000000001",--21919
"001111000110000000110000000000000010",--21920
"001111001110000001000000000000000010",--21921
"111110000110010001000001100000000000",--21922
"001011001010000000110000000000000010",--21923
"011111001101000000100000000000001110",--21924
"001101001000000001000000000000000100",--21925
"001111001010000000110000000000000000",--21926
"001111001010000001000000000000000001",--21927
"001111001010000001010000000000000010",--21928
"001111001000000001100000000000000000",--21929
"111110001100001000110001100000000000",--21930
"001111001000000001100000000000000001",--21931
"111110001100001001000010000000000000",--21932
"111110000110000001000001100000000000",--21933
"001111001000000001000000000000000010",--21934
"111110001000001001010010000000000000",--21935
"111110000110000001000001100000000000",--21936
"001011001010000000110000000000000011",--21937
"000101000000000000000101010111011000",--21938
"010111001101000000100000000000100100",--21939
"001111001010000000110000000000000000",--21940
"001111001010000001000000000000000001",--21941
"001111001010000001010000000000000010",--21942
"111110000110001000110011000000000000",--21943
"001101001000000001110000000000000100",--21944
"001111001110000001110000000000000000",--21945
"111110001100001001110011000000000000",--21946
"111110001000001001000011100000000000",--21947
"001111001110000010000000000000000001",--21948
"111110001110001010000011100000000000",--21949
"111110001100000001110011000000000000",--21950
"111110001010001001010011100000000000",--21951
"001111001110000010000000000000000010",--21952
"111110001110001010000011100000000000",--21953
"111110001100000001110011000000000000",--21954
"001101001000000001110000000000000011",--21955
"011100001111000000000000000000000011",--21956
"101110001101111000000001100000000000",--21957
"011111001101000000110000000000010000",--21958
"000101000000000000000101010111010110",--21959
"111110001000001001010011100000000000",--21960
"001101001000000001000000000000001001",--21961
"001111001000000010000000000000000000",--21962
"111110001110001010000011100000000000",--21963
"111110001100000001110011000000000000",--21964
"111110001010001000110010100000000000",--21965
"001111001000000001110000000000000001",--21966
"111110001010001001110010100000000000",--21967
"111110001100000001010010100000000000",--21968
"111110000110001001000001100000000000",--21969
"001111001000000001000000000000000010",--21970
"111110000110001001000001100000000000",--21971
"111110001010000000110001100000000000",--21972
"011111001101000000110000000000000001",--21973
"111110000110010000010001100000000000",--21974
"001011001010000000110000000000000011",--21975
"101001000100010000100000000000000001",--21976
"010111000101000000000000000010010001",--21977
"001101000100000001000000000101101101",--21978
"001101001000000001010000000000001010",--21979
"001101001000000001100000000000000001",--21980
"001111000110000000110000000000000000",--21981
"001101001000000001110000000000000101",--21982
"001111001110000001000000000000000000",--21983
"111110000110010001000001100000000000",--21984
"001011001010000000110000000000000000",--21985
"001111000110000000110000000000000001",--21986
"001111001110000001000000000000000001",--21987
"111110000110010001000001100000000000",--21988
"001011001010000000110000000000000001",--21989
"001111000110000000110000000000000010",--21990
"001111001110000001000000000000000010",--21991
"111110000110010001000001100000000000",--21992
"001011001010000000110000000000000010",--21993
"011111001101000000100000000000001110",--21994
"001101001000000001000000000000000100",--21995
"001111001010000000110000000000000000",--21996
"001111001010000001000000000000000001",--21997
"001111001010000001010000000000000010",--21998
"001111001000000001100000000000000000",--21999
"111110001100001000110001100000000000",--22000
"001111001000000001100000000000000001",--22001
"111110001100001001000010000000000000",--22002
"111110000110000001000001100000000000",--22003
"001111001000000001000000000000000010",--22004
"111110001000001001010010000000000000",--22005
"111110000110000001000001100000000000",--22006
"001011001010000000110000000000000011",--22007
"000101000000000000000101011000011110",--22008
"010111001101000000100000000000100100",--22009
"001111001010000000110000000000000000",--22010
"001111001010000001000000000000000001",--22011
"001111001010000001010000000000000010",--22012
"111110000110001000110011000000000000",--22013
"001101001000000001110000000000000100",--22014
"001111001110000001110000000000000000",--22015
"111110001100001001110011000000000000",--22016
"111110001000001001000011100000000000",--22017
"001111001110000010000000000000000001",--22018
"111110001110001010000011100000000000",--22019
"111110001100000001110011000000000000",--22020
"111110001010001001010011100000000000",--22021
"001111001110000010000000000000000010",--22022
"111110001110001010000011100000000000",--22023
"111110001100000001110011000000000000",--22024
"001101001000000001110000000000000011",--22025
"011100001111000000000000000000000011",--22026
"101110001101111000000001100000000000",--22027
"011111001101000000110000000000010000",--22028
"000101000000000000000101011000011100",--22029
"111110001000001001010011100000000000",--22030
"001101001000000001000000000000001001",--22031
"001111001000000010000000000000000000",--22032
"111110001110001010000011100000000000",--22033
"111110001100000001110011000000000000",--22034
"111110001010001000110010100000000000",--22035
"001111001000000001110000000000000001",--22036
"111110001010001001110010100000000000",--22037
"111110001100000001010010100000000000",--22038
"111110000110001001000001100000000000",--22039
"001111001000000001000000000000000010",--22040
"111110000110001001000001100000000000",--22041
"111110001010000000110001100000000000",--22042
"011111001101000000110000000000000001",--22043
"111110000110010000010001100000000000",--22044
"001011001010000000110000000000000011",--22045
"101001000100010000100000000000000001",--22046
"010111000101000000000000000001001011",--22047
"001101000100000001000000000101101101",--22048
"001101001000000001010000000000001010",--22049
"001101001000000001100000000000000001",--22050
"001111000110000000110000000000000000",--22051
"001101001000000001110000000000000101",--22052
"001111001110000001000000000000000000",--22053
"111110000110010001000001100000000000",--22054
"001011001010000000110000000000000000",--22055
"001111000110000000110000000000000001",--22056
"001111001110000001000000000000000001",--22057
"111110000110010001000001100000000000",--22058
"001011001010000000110000000000000001",--22059
"001111000110000000110000000000000010",--22060
"001111001110000001000000000000000010",--22061
"111110000110010001000001100000000000",--22062
"001011001010000000110000000000000010",--22063
"011111001101000000100000000000001110",--22064
"001101001000000001000000000000000100",--22065
"001111001010000000110000000000000000",--22066
"001111001010000001000000000000000001",--22067
"001111001010000001010000000000000010",--22068
"001111001000000001100000000000000000",--22069
"111110001100001000110001100000000000",--22070
"001111001000000001100000000000000001",--22071
"111110001100001001000010000000000000",--22072
"111110000110000001000001100000000000",--22073
"001111001000000001000000000000000010",--22074
"111110001000001001010010000000000000",--22075
"111110000110000001000001100000000000",--22076
"001011001010000000110000000000000011",--22077
"000101000000000000000101011001100100",--22078
"010111001101000000100000000000100100",--22079
"001111001010000000110000000000000000",--22080
"001111001010000001000000000000000001",--22081
"001111001010000001010000000000000010",--22082
"111110000110001000110011000000000000",--22083
"001101001000000001110000000000000100",--22084
"001111001110000001110000000000000000",--22085
"111110001100001001110011000000000000",--22086
"111110001000001001000011100000000000",--22087
"001111001110000010000000000000000001",--22088
"111110001110001010000011100000000000",--22089
"111110001100000001110011000000000000",--22090
"111110001010001001010011100000000000",--22091
"001111001110000010000000000000000010",--22092
"111110001110001010000011100000000000",--22093
"111110001100000001110011000000000000",--22094
"001101001000000001110000000000000011",--22095
"011100001111000000000000000000000011",--22096
"101110001101111000000001100000000000",--22097
"011111001101000000110000000000010000",--22098
"000101000000000000000101011001100010",--22099
"111110001000001001010011100000000000",--22100
"001101001000000001000000000000001001",--22101
"001111001000000010000000000000000000",--22102
"111110001110001010000011100000000000",--22103
"111110001100000001110011000000000000",--22104
"111110001010001000110010100000000000",--22105
"001111001000000001110000000000000001",--22106
"111110001010001001110010100000000000",--22107
"111110001100000001010010100000000000",--22108
"111110000110001001000001100000000000",--22109
"001111001000000001000000000000000010",--22110
"111110000110001001000001100000000000",--22111
"111110001010000000110001100000000000",--22112
"011111001101000000110000000000000001",--22113
"111110000110010000010001100000000000",--22114
"001011001010000000110000000000000011",--22115
"101001000100010000100000000000000001",--22116
"101000000111111000000000100000000000",--22117
"001001111100000111111111111111111100",--22118
"101001111100010111100000000000000101",--22119
"000111000000000000000000011001101110",--22120
"101001111100000111100000000000000101",--22121
"001101111100000111111111111111111100",--22122
"101001000000000001000000000001110110",--22123
"001101111100000000011111111111111101",--22124
"001101111100000000100000000000000000",--22125
"001101111100000000111111111111111111",--22126
"000101000000000000000100000011011011",--22127
"001101000010000000110000000000000101",--22128
"001101000010000001000000000000000111",--22129
"001101000010000001010000000000000001",--22130
"001101000010000001100000000000000100",--22131
"001100000110000000100001100000000000",--22132
"001111000110000000110000000000000000",--22133
"001011000000000000110000000100100000",--22134
"001111000110000000110000000000000001",--22135
"001011000000000000110000000100100001",--22136
"001111000110000000110000000000000010",--22137
"001011000000000000110000000100100010",--22138
"001101000010000000010000000000000110",--22139
"001101000010000000010000000000000000",--22140
"001100001000000000100001100000000000",--22141
"001100001010000000100010000000000000",--22142
"001001111100000001100000000000000000",--22143
"001001111100000000101111111111111111",--22144
"001001111100000000111111111111111110",--22145
"001001111100000001001111111111111101",--22146
"001001111100000000011111111111111100",--22147
"010000000011000000000000000011001000",--22148
"001101000000000001010000000011111110",--22149
"001111001000000000110000000000000000",--22150
"001011000000000000110000000100010010",--22151
"001111001000000000110000000000000001",--22152
"001011000000000000110000000100010011",--22153
"001111001000000000110000000000000010",--22154
"001011000000000000110000000100010100",--22155
"001101000000000001110000000110101010",--22156
"101001001110010001110000000000000001",--22157
"001001111100000001011111111111111011",--22158
"010111001111000000000000000010010001",--22159
"001101001110000010000000000101101101",--22160
"001101010000000010010000000000001010",--22161
"001101010000000010100000000000000001",--22162
"001111001000000000110000000000000000",--22163
"001101010000000010110000000000000101",--22164
"001111010110000001000000000000000000",--22165
"111110000110010001000001100000000000",--22166
"001011010010000000110000000000000000",--22167
"001111001000000000110000000000000001",--22168
"001111010110000001000000000000000001",--22169
"111110000110010001000001100000000000",--22170
"001011010010000000110000000000000001",--22171
"001111001000000000110000000000000010",--22172
"001111010110000001000000000000000010",--22173
"111110000110010001000001100000000000",--22174
"001011010010000000110000000000000010",--22175
"011111010101000000100000000000001110",--22176
"001101010000000010000000000000000100",--22177
"001111010010000000110000000000000000",--22178
"001111010010000001000000000000000001",--22179
"001111010010000001010000000000000010",--22180
"001111010000000001100000000000000000",--22181
"111110001100001000110001100000000000",--22182
"001111010000000001100000000000000001",--22183
"111110001100001001000010000000000000",--22184
"111110000110000001000001100000000000",--22185
"001111010000000001000000000000000010",--22186
"111110001000001001010010000000000000",--22187
"111110000110000001000001100000000000",--22188
"001011010010000000110000000000000011",--22189
"000101000000000000000101011011010100",--22190
"010111010101000000100000000000100100",--22191
"001111010010000000110000000000000000",--22192
"001111010010000001000000000000000001",--22193
"001111010010000001010000000000000010",--22194
"111110000110001000110011000000000000",--22195
"001101010000000010110000000000000100",--22196
"001111010110000001110000000000000000",--22197
"111110001100001001110011000000000000",--22198
"111110001000001001000011100000000000",--22199
"001111010110000010000000000000000001",--22200
"111110001110001010000011100000000000",--22201
"111110001100000001110011000000000000",--22202
"111110001010001001010011100000000000",--22203
"001111010110000010000000000000000010",--22204
"111110001110001010000011100000000000",--22205
"111110001100000001110011000000000000",--22206
"001101010000000010110000000000000011",--22207
"011100010111000000000000000000000011",--22208
"101110001101111000000001100000000000",--22209
"011111010101000000110000000000010000",--22210
"000101000000000000000101011011010010",--22211
"111110001000001001010011100000000000",--22212
"001101010000000010000000000000001001",--22213
"001111010000000010000000000000000000",--22214
"111110001110001010000011100000000000",--22215
"111110001100000001110011000000000000",--22216
"111110001010001000110010100000000000",--22217
"001111010000000001110000000000000001",--22218
"111110001010001001110010100000000000",--22219
"111110001100000001010010100000000000",--22220
"111110000110001001000001100000000000",--22221
"001111010000000001000000000000000010",--22222
"111110000110001001000001100000000000",--22223
"111110001010000000110001100000000000",--22224
"011111010101000000110000000000000001",--22225
"111110000110010000010001100000000000",--22226
"001011010010000000110000000000000011",--22227
"101001001110010001110000000000000001",--22228
"010111001111000000000000000001001011",--22229
"001101001110000010000000000101101101",--22230
"001101010000000010010000000000001010",--22231
"001101010000000010100000000000000001",--22232
"001111001000000000110000000000000000",--22233
"001101010000000010110000000000000101",--22234
"001111010110000001000000000000000000",--22235
"111110000110010001000001100000000000",--22236
"001011010010000000110000000000000000",--22237
"001111001000000000110000000000000001",--22238
"001111010110000001000000000000000001",--22239
"111110000110010001000001100000000000",--22240
"001011010010000000110000000000000001",--22241
"001111001000000000110000000000000010",--22242
"001111010110000001000000000000000010",--22243
"111110000110010001000001100000000000",--22244
"001011010010000000110000000000000010",--22245
"011111010101000000100000000000001110",--22246
"001101010000000010000000000000000100",--22247
"001111010010000000110000000000000000",--22248
"001111010010000001000000000000000001",--22249
"001111010010000001010000000000000010",--22250
"001111010000000001100000000000000000",--22251
"111110001100001000110001100000000000",--22252
"001111010000000001100000000000000001",--22253
"111110001100001001000010000000000000",--22254
"111110000110000001000001100000000000",--22255
"001111010000000001000000000000000010",--22256
"111110001000001001010010000000000000",--22257
"111110000110000001000001100000000000",--22258
"001011010010000000110000000000000011",--22259
"000101000000000000000101011100011010",--22260
"010111010101000000100000000000100100",--22261
"001111010010000000110000000000000000",--22262
"001111010010000001000000000000000001",--22263
"001111010010000001010000000000000010",--22264
"111110000110001000110011000000000000",--22265
"001101010000000010110000000000000100",--22266
"001111010110000001110000000000000000",--22267
"111110001100001001110011000000000000",--22268
"111110001000001001000011100000000000",--22269
"001111010110000010000000000000000001",--22270
"111110001110001010000011100000000000",--22271
"111110001100000001110011000000000000",--22272
"111110001010001001010011100000000000",--22273
"001111010110000010000000000000000010",--22274
"111110001110001010000011100000000000",--22275
"111110001100000001110011000000000000",--22276
"001101010000000010110000000000000011",--22277
"011100010111000000000000000000000011",--22278
"101110001101111000000001100000000000",--22279
"011111010101000000110000000000010000",--22280
"000101000000000000000101011100011000",--22281
"111110001000001001010011100000000000",--22282
"001101010000000010000000000000001001",--22283
"001111010000000010000000000000000000",--22284
"111110001110001010000011100000000000",--22285
"111110001100000001110011000000000000",--22286
"111110001010001000110010100000000000",--22287
"001111010000000001110000000000000001",--22288
"111110001010001001110010100000000000",--22289
"111110001100000001010010100000000000",--22290
"111110000110001001000001100000000000",--22291
"001111010000000001000000000000000010",--22292
"111110000110001001000001100000000000",--22293
"111110001010000000110001100000000000",--22294
"011111010101000000110000000000000001",--22295
"111110000110010000010001100000000000",--22296
"001011010010000000110000000000000011",--22297
"101001001110010000100000000000000001",--22298
"101000001001111000000000100000000000",--22299
"001001111100000111111111111111111010",--22300
"101001111100010111100000000000000111",--22301
"000111000000000000000000011001101110",--22302
"101001111100000111100000000000000111",--22303
"001101111100000111111111111111111010",--22304
"001101111100000000011111111111111011",--22305
"001101000010000000100000000001110110",--22306
"001101000100000000100000000000000000",--22307
"001111000100000000110000000000000000",--22308
"001101111100000000111111111111111110",--22309
"001111000110000001000000000000000000",--22310
"111110000110001001000001100000000000",--22311
"001111000100000001000000000000000001",--22312
"001111000110000001010000000000000001",--22313
"111110001000001001010010000000000000",--22314
"111110000110000001000001100000000000",--22315
"001111000100000001000000000000000010",--22316
"001111000110000001010000000000000010",--22317
"111110001000001001010010000000000000",--22318
"111110000110000001000001100000000000",--22319
"011010000111000000000000000000001010",--22320
"001101000010000000010000000001110111",--22321
"101111001001110001001011101111011010",--22322
"101111001001100001000111010000001101",--22323
"111110000110001001000001100000000000",--22324
"001001111100000111111111111111111010",--22325
"101001111100010111100000000000000111",--22326
"000111000000000000000011110001110100",--22327
"101001111100000111100000000000000111",--22328
"001101111100000111111111111111111010",--22329
"000101000000000000000101011101000100",--22330
"001101000010000000010000000001110110",--22331
"101111001001110001000011101111011010",--22332
"101111001001100001000111010000001101",--22333
"111110000110001001000001100000000000",--22334
"001001111100000111111111111111111010",--22335
"101001111100010111100000000000000111",--22336
"000111000000000000000011110001110100",--22337
"101001111100000111100000000000000111",--22338
"001101111100000111111111111111111010",--22339
"101001000000000001000000000001110100",--22340
"001101111100000000011111111111111011",--22341
"001101111100000000101111111111111110",--22342
"001101111100000000111111111111111101",--22343
"001001111100000111111111111111111010",--22344
"101001111100010111100000000000000111",--22345
"000111000000000000000100000011011010",--22346
"101001111100000111100000000000000111",--22347
"001101111100000111111111111111111010",--22348
"001101111100000000011111111111111100",--22349
"010011000011000000010000000011001001",--22350
"001101000000000000100000000011111111",--22351
"001101111100000000111111111111111101",--22352
"001111000110000000110000000000000000",--22353
"001011000000000000110000000100010010",--22354
"001111000110000000110000000000000001",--22355
"001011000000000000110000000100010011",--22356
"001111000110000000110000000000000010",--22357
"001011000000000000110000000100010100",--22358
"001101000000000001000000000110101010",--22359
"101001001000010001000000000000000001",--22360
"001001111100000000101111111111111011",--22361
"010111001001000000000000000010010001",--22362
"001101001000000001010000000101101101",--22363
"001101001010000001100000000000001010",--22364
"001101001010000001110000000000000001",--22365
"001111000110000000110000000000000000",--22366
"001101001010000010000000000000000101",--22367
"001111010000000001000000000000000000",--22368
"111110000110010001000001100000000000",--22369
"001011001100000000110000000000000000",--22370
"001111000110000000110000000000000001",--22371
"001111010000000001000000000000000001",--22372
"111110000110010001000001100000000000",--22373
"001011001100000000110000000000000001",--22374
"001111000110000000110000000000000010",--22375
"001111010000000001000000000000000010",--22376
"111110000110010001000001100000000000",--22377
"001011001100000000110000000000000010",--22378
"011111001111000000100000000000001110",--22379
"001101001010000001010000000000000100",--22380
"001111001100000000110000000000000000",--22381
"001111001100000001000000000000000001",--22382
"001111001100000001010000000000000010",--22383
"001111001010000001100000000000000000",--22384
"111110001100001000110001100000000000",--22385
"001111001010000001100000000000000001",--22386
"111110001100001001000010000000000000",--22387
"111110000110000001000001100000000000",--22388
"001111001010000001000000000000000010",--22389
"111110001000001001010010000000000000",--22390
"111110000110000001000001100000000000",--22391
"001011001100000000110000000000000011",--22392
"000101000000000000000101011110011111",--22393
"010111001111000000100000000000100100",--22394
"001111001100000000110000000000000000",--22395
"001111001100000001000000000000000001",--22396
"001111001100000001010000000000000010",--22397
"111110000110001000110011000000000000",--22398
"001101001010000010000000000000000100",--22399
"001111010000000001110000000000000000",--22400
"111110001100001001110011000000000000",--22401
"111110001000001001000011100000000000",--22402
"001111010000000010000000000000000001",--22403
"111110001110001010000011100000000000",--22404
"111110001100000001110011000000000000",--22405
"111110001010001001010011100000000000",--22406
"001111010000000010000000000000000010",--22407
"111110001110001010000011100000000000",--22408
"111110001100000001110011000000000000",--22409
"001101001010000010000000000000000011",--22410
"011100010001000000000000000000000011",--22411
"101110001101111000000001100000000000",--22412
"011111001111000000110000000000010000",--22413
"000101000000000000000101011110011101",--22414
"111110001000001001010011100000000000",--22415
"001101001010000001010000000000001001",--22416
"001111001010000010000000000000000000",--22417
"111110001110001010000011100000000000",--22418
"111110001100000001110011000000000000",--22419
"111110001010001000110010100000000000",--22420
"001111001010000001110000000000000001",--22421
"111110001010001001110010100000000000",--22422
"111110001100000001010010100000000000",--22423
"111110000110001001000001100000000000",--22424
"001111001010000001000000000000000010",--22425
"111110000110001001000001100000000000",--22426
"111110001010000000110001100000000000",--22427
"011111001111000000110000000000000001",--22428
"111110000110010000010001100000000000",--22429
"001011001100000000110000000000000011",--22430
"101001001000010001000000000000000001",--22431
"010111001001000000000000000001001011",--22432
"001101001000000001010000000101101101",--22433
"001101001010000001100000000000001010",--22434
"001101001010000001110000000000000001",--22435
"001111000110000000110000000000000000",--22436
"001101001010000010000000000000000101",--22437
"001111010000000001000000000000000000",--22438
"111110000110010001000001100000000000",--22439
"001011001100000000110000000000000000",--22440
"001111000110000000110000000000000001",--22441
"001111010000000001000000000000000001",--22442
"111110000110010001000001100000000000",--22443
"001011001100000000110000000000000001",--22444
"001111000110000000110000000000000010",--22445
"001111010000000001000000000000000010",--22446
"111110000110010001000001100000000000",--22447
"001011001100000000110000000000000010",--22448
"011111001111000000100000000000001110",--22449
"001101001010000001010000000000000100",--22450
"001111001100000000110000000000000000",--22451
"001111001100000001000000000000000001",--22452
"001111001100000001010000000000000010",--22453
"001111001010000001100000000000000000",--22454
"111110001100001000110001100000000000",--22455
"001111001010000001100000000000000001",--22456
"111110001100001001000010000000000000",--22457
"111110000110000001000001100000000000",--22458
"001111001010000001000000000000000010",--22459
"111110001000001001010010000000000000",--22460
"111110000110000001000001100000000000",--22461
"001011001100000000110000000000000011",--22462
"000101000000000000000101011111100101",--22463
"010111001111000000100000000000100100",--22464
"001111001100000000110000000000000000",--22465
"001111001100000001000000000000000001",--22466
"001111001100000001010000000000000010",--22467
"111110000110001000110011000000000000",--22468
"001101001010000010000000000000000100",--22469
"001111010000000001110000000000000000",--22470
"111110001100001001110011000000000000",--22471
"111110001000001001000011100000000000",--22472
"001111010000000010000000000000000001",--22473
"111110001110001010000011100000000000",--22474
"111110001100000001110011000000000000",--22475
"111110001010001001010011100000000000",--22476
"001111010000000010000000000000000010",--22477
"111110001110001010000011100000000000",--22478
"111110001100000001110011000000000000",--22479
"001101001010000010000000000000000011",--22480
"011100010001000000000000000000000011",--22481
"101110001101111000000001100000000000",--22482
"011111001111000000110000000000010000",--22483
"000101000000000000000101011111100011",--22484
"111110001000001001010011100000000000",--22485
"001101001010000001010000000000001001",--22486
"001111001010000010000000000000000000",--22487
"111110001110001010000011100000000000",--22488
"111110001100000001110011000000000000",--22489
"111110001010001000110010100000000000",--22490
"001111001010000001110000000000000001",--22491
"111110001010001001110010100000000000",--22492
"111110001100000001010010100000000000",--22493
"111110000110001001000001100000000000",--22494
"001111001010000001000000000000000010",--22495
"111110000110001001000001100000000000",--22496
"111110001010000000110001100000000000",--22497
"011111001111000000110000000000000001",--22498
"111110000110010000010001100000000000",--22499
"001011001100000000110000000000000011",--22500
"101001001000010000100000000000000001",--22501
"101000000111111000000000100000000000",--22502
"001001111100000111111111111111111010",--22503
"101001111100010111100000000000000111",--22504
"000111000000000000000000011001101110",--22505
"101001111100000111100000000000000111",--22506
"001101111100000111111111111111111010",--22507
"001101111100000000011111111111111011",--22508
"001101000010000000100000000001110110",--22509
"001101000100000000100000000000000000",--22510
"001111000100000000110000000000000000",--22511
"001101111100000000111111111111111110",--22512
"001111000110000001000000000000000000",--22513
"111110000110001001000001100000000000",--22514
"001111000100000001000000000000000001",--22515
"001111000110000001010000000000000001",--22516
"111110001000001001010010000000000000",--22517
"111110000110000001000001100000000000",--22518
"001111000100000001000000000000000010",--22519
"001111000110000001010000000000000010",--22520
"111110001000001001010010000000000000",--22521
"111110000110000001000001100000000000",--22522
"011010000111000000000000000000001010",--22523
"001101000010000000010000000001110111",--22524
"101111001001110001001011101111011010",--22525
"101111001001100001000111010000001101",--22526
"111110000110001001000001100000000000",--22527
"001001111100000111111111111111111010",--22528
"101001111100010111100000000000000111",--22529
"000111000000000000000011110001110100",--22530
"101001111100000111100000000000000111",--22531
"001101111100000111111111111111111010",--22532
"000101000000000000000101100000001111",--22533
"001101000010000000010000000001110110",--22534
"101111001001110001000011101111011010",--22535
"101111001001100001000111010000001101",--22536
"111110000110001001000001100000000000",--22537
"001001111100000111111111111111111010",--22538
"101001111100010111100000000000000111",--22539
"000111000000000000000011110001110100",--22540
"101001111100000111100000000000000111",--22541
"001101111100000111111111111111111010",--22542
"101001000000000001000000000001110100",--22543
"001101111100000000011111111111111011",--22544
"001101111100000000101111111111111110",--22545
"001101111100000000111111111111111101",--22546
"001001111100000111111111111111111010",--22547
"101001111100010111100000000000000111",--22548
"000111000000000000000100000011011010",--22549
"101001111100000111100000000000000111",--22550
"001101111100000111111111111111111010",--22551
"001101111100000000011111111111111100",--22552
"010011000011000000100000000011001001",--22553
"001101000000000000100000000100000000",--22554
"001101111100000000111111111111111101",--22555
"001111000110000000110000000000000000",--22556
"001011000000000000110000000100010010",--22557
"001111000110000000110000000000000001",--22558
"001011000000000000110000000100010011",--22559
"001111000110000000110000000000000010",--22560
"001011000000000000110000000100010100",--22561
"001101000000000001000000000110101010",--22562
"101001001000010001000000000000000001",--22563
"001001111100000000101111111111111011",--22564
"010111001001000000000000000010010001",--22565
"001101001000000001010000000101101101",--22566
"001101001010000001100000000000001010",--22567
"001101001010000001110000000000000001",--22568
"001111000110000000110000000000000000",--22569
"001101001010000010000000000000000101",--22570
"001111010000000001000000000000000000",--22571
"111110000110010001000001100000000000",--22572
"001011001100000000110000000000000000",--22573
"001111000110000000110000000000000001",--22574
"001111010000000001000000000000000001",--22575
"111110000110010001000001100000000000",--22576
"001011001100000000110000000000000001",--22577
"001111000110000000110000000000000010",--22578
"001111010000000001000000000000000010",--22579
"111110000110010001000001100000000000",--22580
"001011001100000000110000000000000010",--22581
"011111001111000000100000000000001110",--22582
"001101001010000001010000000000000100",--22583
"001111001100000000110000000000000000",--22584
"001111001100000001000000000000000001",--22585
"001111001100000001010000000000000010",--22586
"001111001010000001100000000000000000",--22587
"111110001100001000110001100000000000",--22588
"001111001010000001100000000000000001",--22589
"111110001100001001000010000000000000",--22590
"111110000110000001000001100000000000",--22591
"001111001010000001000000000000000010",--22592
"111110001000001001010010000000000000",--22593
"111110000110000001000001100000000000",--22594
"001011001100000000110000000000000011",--22595
"000101000000000000000101100001101010",--22596
"010111001111000000100000000000100100",--22597
"001111001100000000110000000000000000",--22598
"001111001100000001000000000000000001",--22599
"001111001100000001010000000000000010",--22600
"111110000110001000110011000000000000",--22601
"001101001010000010000000000000000100",--22602
"001111010000000001110000000000000000",--22603
"111110001100001001110011000000000000",--22604
"111110001000001001000011100000000000",--22605
"001111010000000010000000000000000001",--22606
"111110001110001010000011100000000000",--22607
"111110001100000001110011000000000000",--22608
"111110001010001001010011100000000000",--22609
"001111010000000010000000000000000010",--22610
"111110001110001010000011100000000000",--22611
"111110001100000001110011000000000000",--22612
"001101001010000010000000000000000011",--22613
"011100010001000000000000000000000011",--22614
"101110001101111000000001100000000000",--22615
"011111001111000000110000000000010000",--22616
"000101000000000000000101100001101000",--22617
"111110001000001001010011100000000000",--22618
"001101001010000001010000000000001001",--22619
"001111001010000010000000000000000000",--22620
"111110001110001010000011100000000000",--22621
"111110001100000001110011000000000000",--22622
"111110001010001000110010100000000000",--22623
"001111001010000001110000000000000001",--22624
"111110001010001001110010100000000000",--22625
"111110001100000001010010100000000000",--22626
"111110000110001001000001100000000000",--22627
"001111001010000001000000000000000010",--22628
"111110000110001001000001100000000000",--22629
"111110001010000000110001100000000000",--22630
"011111001111000000110000000000000001",--22631
"111110000110010000010001100000000000",--22632
"001011001100000000110000000000000011",--22633
"101001001000010001000000000000000001",--22634
"010111001001000000000000000001001011",--22635
"001101001000000001010000000101101101",--22636
"001101001010000001100000000000001010",--22637
"001101001010000001110000000000000001",--22638
"001111000110000000110000000000000000",--22639
"001101001010000010000000000000000101",--22640
"001111010000000001000000000000000000",--22641
"111110000110010001000001100000000000",--22642
"001011001100000000110000000000000000",--22643
"001111000110000000110000000000000001",--22644
"001111010000000001000000000000000001",--22645
"111110000110010001000001100000000000",--22646
"001011001100000000110000000000000001",--22647
"001111000110000000110000000000000010",--22648
"001111010000000001000000000000000010",--22649
"111110000110010001000001100000000000",--22650
"001011001100000000110000000000000010",--22651
"011111001111000000100000000000001110",--22652
"001101001010000001010000000000000100",--22653
"001111001100000000110000000000000000",--22654
"001111001100000001000000000000000001",--22655
"001111001100000001010000000000000010",--22656
"001111001010000001100000000000000000",--22657
"111110001100001000110001100000000000",--22658
"001111001010000001100000000000000001",--22659
"111110001100001001000010000000000000",--22660
"111110000110000001000001100000000000",--22661
"001111001010000001000000000000000010",--22662
"111110001000001001010010000000000000",--22663
"111110000110000001000001100000000000",--22664
"001011001100000000110000000000000011",--22665
"000101000000000000000101100010110000",--22666
"010111001111000000100000000000100100",--22667
"001111001100000000110000000000000000",--22668
"001111001100000001000000000000000001",--22669
"001111001100000001010000000000000010",--22670
"111110000110001000110011000000000000",--22671
"001101001010000010000000000000000100",--22672
"001111010000000001110000000000000000",--22673
"111110001100001001110011000000000000",--22674
"111110001000001001000011100000000000",--22675
"001111010000000010000000000000000001",--22676
"111110001110001010000011100000000000",--22677
"111110001100000001110011000000000000",--22678
"111110001010001001010011100000000000",--22679
"001111010000000010000000000000000010",--22680
"111110001110001010000011100000000000",--22681
"111110001100000001110011000000000000",--22682
"001101001010000010000000000000000011",--22683
"011100010001000000000000000000000011",--22684
"101110001101111000000001100000000000",--22685
"011111001111000000110000000000010000",--22686
"000101000000000000000101100010101110",--22687
"111110001000001001010011100000000000",--22688
"001101001010000001010000000000001001",--22689
"001111001010000010000000000000000000",--22690
"111110001110001010000011100000000000",--22691
"111110001100000001110011000000000000",--22692
"111110001010001000110010100000000000",--22693
"001111001010000001110000000000000001",--22694
"111110001010001001110010100000000000",--22695
"111110001100000001010010100000000000",--22696
"111110000110001001000001100000000000",--22697
"001111001010000001000000000000000010",--22698
"111110000110001001000001100000000000",--22699
"111110001010000000110001100000000000",--22700
"011111001111000000110000000000000001",--22701
"111110000110010000010001100000000000",--22702
"001011001100000000110000000000000011",--22703
"101001001000010000100000000000000001",--22704
"101000000111111000000000100000000000",--22705
"001001111100000111111111111111111010",--22706
"101001111100010111100000000000000111",--22707
"000111000000000000000000011001101110",--22708
"101001111100000111100000000000000111",--22709
"001101111100000111111111111111111010",--22710
"001101111100000000011111111111111011",--22711
"001101000010000000100000000001110110",--22712
"001101000100000000100000000000000000",--22713
"001111000100000000110000000000000000",--22714
"001101111100000000111111111111111110",--22715
"001111000110000001000000000000000000",--22716
"111110000110001001000001100000000000",--22717
"001111000100000001000000000000000001",--22718
"001111000110000001010000000000000001",--22719
"111110001000001001010010000000000000",--22720
"111110000110000001000001100000000000",--22721
"001111000100000001000000000000000010",--22722
"001111000110000001010000000000000010",--22723
"111110001000001001010010000000000000",--22724
"111110000110000001000001100000000000",--22725
"011010000111000000000000000000001010",--22726
"001101000010000000010000000001110111",--22727
"101111001001110001001011101111011010",--22728
"101111001001100001000111010000001101",--22729
"111110000110001001000001100000000000",--22730
"001001111100000111111111111111111010",--22731
"101001111100010111100000000000000111",--22732
"000111000000000000000011110001110100",--22733
"101001111100000111100000000000000111",--22734
"001101111100000111111111111111111010",--22735
"000101000000000000000101100011011010",--22736
"001101000010000000010000000001110110",--22737
"101111001001110001000011101111011010",--22738
"101111001001100001000111010000001101",--22739
"111110000110001001000001100000000000",--22740
"001001111100000111111111111111111010",--22741
"101001111100010111100000000000000111",--22742
"000111000000000000000011110001110100",--22743
"101001111100000111100000000000000111",--22744
"001101111100000111111111111111111010",--22745
"101001000000000001000000000001110100",--22746
"001101111100000000011111111111111011",--22747
"001101111100000000101111111111111110",--22748
"001101111100000000111111111111111101",--22749
"001001111100000111111111111111111010",--22750
"101001111100010111100000000000000111",--22751
"000111000000000000000100000011011010",--22752
"101001111100000111100000000000000111",--22753
"001101111100000111111111111111111010",--22754
"001101111100000000011111111111111100",--22755
"010011000011000000110000000011001001",--22756
"001101000000000000100000000100000001",--22757
"001101111100000000111111111111111101",--22758
"001111000110000000110000000000000000",--22759
"001011000000000000110000000100010010",--22760
"001111000110000000110000000000000001",--22761
"001011000000000000110000000100010011",--22762
"001111000110000000110000000000000010",--22763
"001011000000000000110000000100010100",--22764
"001101000000000001000000000110101010",--22765
"101001001000010001000000000000000001",--22766
"001001111100000000101111111111111011",--22767
"010111001001000000000000000010010001",--22768
"001101001000000001010000000101101101",--22769
"001101001010000001100000000000001010",--22770
"001101001010000001110000000000000001",--22771
"001111000110000000110000000000000000",--22772
"001101001010000010000000000000000101",--22773
"001111010000000001000000000000000000",--22774
"111110000110010001000001100000000000",--22775
"001011001100000000110000000000000000",--22776
"001111000110000000110000000000000001",--22777
"001111010000000001000000000000000001",--22778
"111110000110010001000001100000000000",--22779
"001011001100000000110000000000000001",--22780
"001111000110000000110000000000000010",--22781
"001111010000000001000000000000000010",--22782
"111110000110010001000001100000000000",--22783
"001011001100000000110000000000000010",--22784
"011111001111000000100000000000001110",--22785
"001101001010000001010000000000000100",--22786
"001111001100000000110000000000000000",--22787
"001111001100000001000000000000000001",--22788
"001111001100000001010000000000000010",--22789
"001111001010000001100000000000000000",--22790
"111110001100001000110001100000000000",--22791
"001111001010000001100000000000000001",--22792
"111110001100001001000010000000000000",--22793
"111110000110000001000001100000000000",--22794
"001111001010000001000000000000000010",--22795
"111110001000001001010010000000000000",--22796
"111110000110000001000001100000000000",--22797
"001011001100000000110000000000000011",--22798
"000101000000000000000101100100110101",--22799
"010111001111000000100000000000100100",--22800
"001111001100000000110000000000000000",--22801
"001111001100000001000000000000000001",--22802
"001111001100000001010000000000000010",--22803
"111110000110001000110011000000000000",--22804
"001101001010000010000000000000000100",--22805
"001111010000000001110000000000000000",--22806
"111110001100001001110011000000000000",--22807
"111110001000001001000011100000000000",--22808
"001111010000000010000000000000000001",--22809
"111110001110001010000011100000000000",--22810
"111110001100000001110011000000000000",--22811
"111110001010001001010011100000000000",--22812
"001111010000000010000000000000000010",--22813
"111110001110001010000011100000000000",--22814
"111110001100000001110011000000000000",--22815
"001101001010000010000000000000000011",--22816
"011100010001000000000000000000000011",--22817
"101110001101111000000001100000000000",--22818
"011111001111000000110000000000010000",--22819
"000101000000000000000101100100110011",--22820
"111110001000001001010011100000000000",--22821
"001101001010000001010000000000001001",--22822
"001111001010000010000000000000000000",--22823
"111110001110001010000011100000000000",--22824
"111110001100000001110011000000000000",--22825
"111110001010001000110010100000000000",--22826
"001111001010000001110000000000000001",--22827
"111110001010001001110010100000000000",--22828
"111110001100000001010010100000000000",--22829
"111110000110001001000001100000000000",--22830
"001111001010000001000000000000000010",--22831
"111110000110001001000001100000000000",--22832
"111110001010000000110001100000000000",--22833
"011111001111000000110000000000000001",--22834
"111110000110010000010001100000000000",--22835
"001011001100000000110000000000000011",--22836
"101001001000010001000000000000000001",--22837
"010111001001000000000000000001001011",--22838
"001101001000000001010000000101101101",--22839
"001101001010000001100000000000001010",--22840
"001101001010000001110000000000000001",--22841
"001111000110000000110000000000000000",--22842
"001101001010000010000000000000000101",--22843
"001111010000000001000000000000000000",--22844
"111110000110010001000001100000000000",--22845
"001011001100000000110000000000000000",--22846
"001111000110000000110000000000000001",--22847
"001111010000000001000000000000000001",--22848
"111110000110010001000001100000000000",--22849
"001011001100000000110000000000000001",--22850
"001111000110000000110000000000000010",--22851
"001111010000000001000000000000000010",--22852
"111110000110010001000001100000000000",--22853
"001011001100000000110000000000000010",--22854
"011111001111000000100000000000001110",--22855
"001101001010000001010000000000000100",--22856
"001111001100000000110000000000000000",--22857
"001111001100000001000000000000000001",--22858
"001111001100000001010000000000000010",--22859
"001111001010000001100000000000000000",--22860
"111110001100001000110001100000000000",--22861
"001111001010000001100000000000000001",--22862
"111110001100001001000010000000000000",--22863
"111110000110000001000001100000000000",--22864
"001111001010000001000000000000000010",--22865
"111110001000001001010010000000000000",--22866
"111110000110000001000001100000000000",--22867
"001011001100000000110000000000000011",--22868
"000101000000000000000101100101111011",--22869
"010111001111000000100000000000100100",--22870
"001111001100000000110000000000000000",--22871
"001111001100000001000000000000000001",--22872
"001111001100000001010000000000000010",--22873
"111110000110001000110011000000000000",--22874
"001101001010000010000000000000000100",--22875
"001111010000000001110000000000000000",--22876
"111110001100001001110011000000000000",--22877
"111110001000001001000011100000000000",--22878
"001111010000000010000000000000000001",--22879
"111110001110001010000011100000000000",--22880
"111110001100000001110011000000000000",--22881
"111110001010001001010011100000000000",--22882
"001111010000000010000000000000000010",--22883
"111110001110001010000011100000000000",--22884
"111110001100000001110011000000000000",--22885
"001101001010000010000000000000000011",--22886
"011100010001000000000000000000000011",--22887
"101110001101111000000001100000000000",--22888
"011111001111000000110000000000010000",--22889
"000101000000000000000101100101111001",--22890
"111110001000001001010011100000000000",--22891
"001101001010000001010000000000001001",--22892
"001111001010000010000000000000000000",--22893
"111110001110001010000011100000000000",--22894
"111110001100000001110011000000000000",--22895
"111110001010001000110010100000000000",--22896
"001111001010000001110000000000000001",--22897
"111110001010001001110010100000000000",--22898
"111110001100000001010010100000000000",--22899
"111110000110001001000001100000000000",--22900
"001111001010000001000000000000000010",--22901
"111110000110001001000001100000000000",--22902
"111110001010000000110001100000000000",--22903
"011111001111000000110000000000000001",--22904
"111110000110010000010001100000000000",--22905
"001011001100000000110000000000000011",--22906
"101001001000010000100000000000000001",--22907
"101000000111111000000000100000000000",--22908
"001001111100000111111111111111111010",--22909
"101001111100010111100000000000000111",--22910
"000111000000000000000000011001101110",--22911
"101001111100000111100000000000000111",--22912
"001101111100000111111111111111111010",--22913
"001101111100000000011111111111111011",--22914
"001101000010000000100000000001110110",--22915
"001101000100000000100000000000000000",--22916
"001111000100000000110000000000000000",--22917
"001101111100000000111111111111111110",--22918
"001111000110000001000000000000000000",--22919
"111110000110001001000001100000000000",--22920
"001111000100000001000000000000000001",--22921
"001111000110000001010000000000000001",--22922
"111110001000001001010010000000000000",--22923
"111110000110000001000001100000000000",--22924
"001111000100000001000000000000000010",--22925
"001111000110000001010000000000000010",--22926
"111110001000001001010010000000000000",--22927
"111110000110000001000001100000000000",--22928
"011010000111000000000000000000001010",--22929
"001101000010000000010000000001110111",--22930
"101111001001110001001011101111011010",--22931
"101111001001100001000111010000001101",--22932
"111110000110001001000001100000000000",--22933
"001001111100000111111111111111111010",--22934
"101001111100010111100000000000000111",--22935
"000111000000000000000011110001110100",--22936
"101001111100000111100000000000000111",--22937
"001101111100000111111111111111111010",--22938
"000101000000000000000101100110100101",--22939
"001101000010000000010000000001110110",--22940
"101111001001110001000011101111011010",--22941
"101111001001100001000111010000001101",--22942
"111110000110001001000001100000000000",--22943
"001001111100000111111111111111111010",--22944
"101001111100010111100000000000000111",--22945
"000111000000000000000011110001110100",--22946
"101001111100000111100000000000000111",--22947
"001101111100000111111111111111111010",--22948
"101001000000000001000000000001110100",--22949
"001101111100000000011111111111111011",--22950
"001101111100000000101111111111111110",--22951
"001101111100000000111111111111111101",--22952
"001001111100000111111111111111111010",--22953
"101001111100010111100000000000000111",--22954
"000111000000000000000100000011011010",--22955
"101001111100000111100000000000000111",--22956
"001101111100000111111111111111111010",--22957
"001101111100000000011111111111111100",--22958
"010011000011000001000000000011001010",--22959
"001101000000000000010000000100000010",--22960
"001101111100000000101111111111111101",--22961
"001111000100000000110000000000000000",--22962
"001011000000000000110000000100010010",--22963
"001111000100000000110000000000000001",--22964
"001011000000000000110000000100010011",--22965
"001111000100000000110000000000000010",--22966
"001011000000000000110000000100010100",--22967
"001101000000000000110000000110101010",--22968
"101001000110010000110000000000000001",--22969
"001001111100000000011111111111111011",--22970
"010111000111000000000000000010010010",--22971
"001101000110000001000000000101101101",--22972
"001101001000000001010000000000001010",--22973
"001101001000000001100000000000000001",--22974
"001111000100000000110000000000000000",--22975
"001101001000000001110000000000000101",--22976
"001111001110000001000000000000000000",--22977
"111110000110010001000001100000000000",--22978
"001011001010000000110000000000000000",--22979
"001111000100000000110000000000000001",--22980
"001111001110000001000000000000000001",--22981
"111110000110010001000001100000000000",--22982
"001011001010000000110000000000000001",--22983
"001111000100000000110000000000000010",--22984
"001111001110000001000000000000000010",--22985
"111110000110010001000001100000000000",--22986
"001011001010000000110000000000000010",--22987
"011111001101000000100000000000001110",--22988
"001101001000000001000000000000000100",--22989
"001111001010000000110000000000000000",--22990
"001111001010000001000000000000000001",--22991
"001111001010000001010000000000000010",--22992
"001111001000000001100000000000000000",--22993
"111110001100001000110001100000000000",--22994
"001111001000000001100000000000000001",--22995
"111110001100001001000010000000000000",--22996
"111110000110000001000001100000000000",--22997
"001111001000000001000000000000000010",--22998
"111110001000001001010010000000000000",--22999
"111110000110000001000001100000000000",--23000
"001011001010000000110000000000000011",--23001
"000101000000000000000101101000000000",--23002
"010111001101000000100000000000100100",--23003
"001111001010000000110000000000000000",--23004
"001111001010000001000000000000000001",--23005
"001111001010000001010000000000000010",--23006
"111110000110001000110011000000000000",--23007
"001101001000000001110000000000000100",--23008
"001111001110000001110000000000000000",--23009
"111110001100001001110011000000000000",--23010
"111110001000001001000011100000000000",--23011
"001111001110000010000000000000000001",--23012
"111110001110001010000011100000000000",--23013
"111110001100000001110011000000000000",--23014
"111110001010001001010011100000000000",--23015
"001111001110000010000000000000000010",--23016
"111110001110001010000011100000000000",--23017
"111110001100000001110011000000000000",--23018
"001101001000000001110000000000000011",--23019
"011100001111000000000000000000000011",--23020
"101110001101111000000001100000000000",--23021
"011111001101000000110000000000010000",--23022
"000101000000000000000101100111111110",--23023
"111110001000001001010011100000000000",--23024
"001101001000000001000000000000001001",--23025
"001111001000000010000000000000000000",--23026
"111110001110001010000011100000000000",--23027
"111110001100000001110011000000000000",--23028
"111110001010001000110010100000000000",--23029
"001111001000000001110000000000000001",--23030
"111110001010001001110010100000000000",--23031
"111110001100000001010010100000000000",--23032
"111110000110001001000001100000000000",--23033
"001111001000000001000000000000000010",--23034
"111110000110001001000001100000000000",--23035
"111110001010000000110001100000000000",--23036
"011111001101000000110000000000000001",--23037
"111110000110010000010001100000000000",--23038
"001011001010000000110000000000000011",--23039
"101001000110010000110000000000000001",--23040
"010111000111000000000000000001001100",--23041
"001101000110000001000000000101101101",--23042
"001101001000000001010000000000001010",--23043
"001101001000000001100000000000000001",--23044
"001111000100000000110000000000000000",--23045
"001101001000000001110000000000000101",--23046
"001111001110000001000000000000000000",--23047
"111110000110010001000001100000000000",--23048
"001011001010000000110000000000000000",--23049
"001111000100000000110000000000000001",--23050
"001111001110000001000000000000000001",--23051
"111110000110010001000001100000000000",--23052
"001011001010000000110000000000000001",--23053
"001111000100000000110000000000000010",--23054
"001111001110000001000000000000000010",--23055
"111110000110010001000001100000000000",--23056
"001011001010000000110000000000000010",--23057
"011111001101000000100000000000001110",--23058
"001101001000000001000000000000000100",--23059
"001111001010000000110000000000000000",--23060
"001111001010000001000000000000000001",--23061
"001111001010000001010000000000000010",--23062
"001111001000000001100000000000000000",--23063
"111110001100001000110001100000000000",--23064
"001111001000000001100000000000000001",--23065
"111110001100001001000010000000000000",--23066
"111110000110000001000001100000000000",--23067
"001111001000000001000000000000000010",--23068
"111110001000001001010010000000000000",--23069
"111110000110000001000001100000000000",--23070
"001011001010000000110000000000000011",--23071
"000101000000000000000101101001000110",--23072
"010111001101000000100000000000100100",--23073
"001111001010000000110000000000000000",--23074
"001111001010000001000000000000000001",--23075
"001111001010000001010000000000000010",--23076
"111110000110001000110011000000000000",--23077
"001101001000000001110000000000000100",--23078
"001111001110000001110000000000000000",--23079
"111110001100001001110011000000000000",--23080
"111110001000001001000011100000000000",--23081
"001111001110000010000000000000000001",--23082
"111110001110001010000011100000000000",--23083
"111110001100000001110011000000000000",--23084
"111110001010001001010011100000000000",--23085
"001111001110000010000000000000000010",--23086
"111110001110001010000011100000000000",--23087
"111110001100000001110011000000000000",--23088
"001101001000000001110000000000000011",--23089
"011100001111000000000000000000000011",--23090
"101110001101111000000001100000000000",--23091
"011111001101000000110000000000010000",--23092
"000101000000000000000101101001000100",--23093
"111110001000001001010011100000000000",--23094
"001101001000000001000000000000001001",--23095
"001111001000000010000000000000000000",--23096
"111110001110001010000011100000000000",--23097
"111110001100000001110011000000000000",--23098
"111110001010001000110010100000000000",--23099
"001111001000000001110000000000000001",--23100
"111110001010001001110010100000000000",--23101
"111110001100000001010010100000000000",--23102
"111110000110001001000001100000000000",--23103
"001111001000000001000000000000000010",--23104
"111110000110001001000001100000000000",--23105
"111110001010000000110001100000000000",--23106
"011111001101000000110000000000000001",--23107
"111110000110010000010001100000000000",--23108
"001011001010000000110000000000000011",--23109
"101001000110010000110000000000000001",--23110
"101000000101111000000000100000000000",--23111
"101000000111111000000001000000000000",--23112
"001001111100000111111111111111111010",--23113
"101001111100010111100000000000000111",--23114
"000111000000000000000000011001101110",--23115
"101001111100000111100000000000000111",--23116
"001101111100000111111111111111111010",--23117
"001101111100000000011111111111111011",--23118
"001101000010000000100000000001110110",--23119
"001101000100000000100000000000000000",--23120
"001111000100000000110000000000000000",--23121
"001101111100000000111111111111111110",--23122
"001111000110000001000000000000000000",--23123
"111110000110001001000001100000000000",--23124
"001111000100000001000000000000000001",--23125
"001111000110000001010000000000000001",--23126
"111110001000001001010010000000000000",--23127
"111110000110000001000001100000000000",--23128
"001111000100000001000000000000000010",--23129
"001111000110000001010000000000000010",--23130
"111110001000001001010010000000000000",--23131
"111110000110000001000001100000000000",--23132
"011010000111000000000000000000001010",--23133
"001101000010000000010000000001110111",--23134
"101111001001110001001011101111011010",--23135
"101111001001100001000111010000001101",--23136
"111110000110001001000001100000000000",--23137
"001001111100000111111111111111111010",--23138
"101001111100010111100000000000000111",--23139
"000111000000000000000011110001110100",--23140
"101001111100000111100000000000000111",--23141
"001101111100000111111111111111111010",--23142
"000101000000000000000101101001110001",--23143
"001101000010000000010000000001110110",--23144
"101111001001110001000011101111011010",--23145
"101111001001100001000111010000001101",--23146
"111110000110001001000001100000000000",--23147
"001001111100000111111111111111111010",--23148
"101001111100010111100000000000000111",--23149
"000111000000000000000011110001110100",--23150
"101001111100000111100000000000000111",--23151
"001101111100000111111111111111111010",--23152
"101001000000000001000000000001110100",--23153
"001101111100000000011111111111111011",--23154
"001101111100000000101111111111111110",--23155
"001101111100000000111111111111111101",--23156
"001001111100000111111111111111111010",--23157
"101001111100010111100000000000000111",--23158
"000111000000000000000100000011011010",--23159
"101001111100000111100000000000000111",--23160
"001101111100000111111111111111111010",--23161
"001101111100000000011111111111111111",--23162
"001101111100000000100000000000000000",--23163
"001100000100000000010000100000000000",--23164
"001111000000000000110000000100011101",--23165
"001111000010000001000000000000000000",--23166
"001111000000000001010000000100100000",--23167
"111110001000001001010010000000000000",--23168
"111110000110000001000001100000000000",--23169
"001011000000000000110000000100011101",--23170
"001111000000000000110000000100011110",--23171
"001111000010000001000000000000000001",--23172
"001111000000000001010000000100100001",--23173
"111110001000001001010010000000000000",--23174
"111110000110000001000001100000000000",--23175
"001011000000000000110000000100011110",--23176
"001111000000000000110000000100011111",--23177
"001111000010000001000000000000000010",--23178
"001111000000000001010000000100100010",--23179
"111110001000001001010010000000000000",--23180
"111110000110000001000001100000000000",--23181
"001011000000000000110000000100011111",--23182
"000100000000000000001111100000000000",--23183
"011011000100000001011111100000000000",--23184
"001101000010000000110000000000000010",--23185
"001100000110000000100010000000000000",--23186
"010111001000000000001111100000000000",--23187
"001101000010000001000000000000000011",--23188
"001100001000000000100010100000000000",--23189
"001001111100000000010000000000000000",--23190
"001001111100000001001111111111111111",--23191
"001001111100000000111111111111111110",--23192
"001001111100000000101111111111111101",--23193
"010000001011000000000000010011001100",--23194
"001101000010000001010000000000000101",--23195
"001101000010000001100000000000000111",--23196
"001101000010000001110000000000000001",--23197
"001101000010000010000000000000000100",--23198
"001100001010000000100010100000000000",--23199
"001111001010000000110000000000000000",--23200
"001011000000000000110000000100100000",--23201
"001111001010000000110000000000000001",--23202
"001011000000000000110000000100100001",--23203
"001111001010000000110000000000000010",--23204
"001011000000000000110000000100100010",--23205
"001101000010000001010000000000000110",--23206
"001101001010000001010000000000000000",--23207
"001100001100000000100011000000000000",--23208
"001100001110000000100011100000000000",--23209
"001001111100000010001111111111111100",--23210
"001001111100000001101111111111111011",--23211
"001001111100000001111111111111111010",--23212
"001001111100000001011111111111111001",--23213
"010000001011000000000000000011101011",--23214
"001101000000000010010000000011111110",--23215
"001111001110000000110000000000000000",--23216
"001011000000000000110000000100010010",--23217
"001111001110000000110000000000000001",--23218
"001011000000000000110000000100010011",--23219
"001111001110000000110000000000000010",--23220
"001011000000000000110000000100010100",--23221
"001101000000000010100000000110101010",--23222
"101001010100010010100000000000000001",--23223
"001001111100000010011111111111111000",--23224
"010111010101000000000000000011010111",--23225
"001101010100000010110000000101101101",--23226
"001101010110000011000000000000001010",--23227
"001101010110000011010000000000000001",--23228
"001111001110000000110000000000000000",--23229
"001101010110000011100000000000000101",--23230
"001111011100000001000000000000000000",--23231
"111110000110010001000001100000000000",--23232
"001011011000000000110000000000000000",--23233
"001111001110000000110000000000000001",--23234
"001111011100000001000000000000000001",--23235
"111110000110010001000001100000000000",--23236
"001011011000000000110000000000000001",--23237
"001111001110000000110000000000000010",--23238
"001111011100000001000000000000000010",--23239
"111110000110010001000001100000000000",--23240
"001011011000000000110000000000000010",--23241
"011111011011000000100000000000001110",--23242
"001101010110000010110000000000000100",--23243
"001111011000000000110000000000000000",--23244
"001111011000000001000000000000000001",--23245
"001111011000000001010000000000000010",--23246
"001111010110000001100000000000000000",--23247
"111110001100001000110001100000000000",--23248
"001111010110000001100000000000000001",--23249
"111110001100001001000010000000000000",--23250
"111110000110000001000001100000000000",--23251
"001111010110000001000000000000000010",--23252
"111110001000001001010010000000000000",--23253
"111110000110000001000001100000000000",--23254
"001011011000000000110000000000000011",--23255
"000101000000000000000101101011111110",--23256
"010111011011000000100000000000100100",--23257
"001111011000000000110000000000000000",--23258
"001111011000000001000000000000000001",--23259
"001111011000000001010000000000000010",--23260
"111110000110001000110011000000000000",--23261
"001101010110000011100000000000000100",--23262
"001111011100000001110000000000000000",--23263
"111110001100001001110011000000000000",--23264
"111110001000001001000011100000000000",--23265
"001111011100000010000000000000000001",--23266
"111110001110001010000011100000000000",--23267
"111110001100000001110011000000000000",--23268
"111110001010001001010011100000000000",--23269
"001111011100000010000000000000000010",--23270
"111110001110001010000011100000000000",--23271
"111110001100000001110011000000000000",--23272
"001101010110000011100000000000000011",--23273
"011100011101000000000000000000000011",--23274
"101110001101111000000001100000000000",--23275
"011111011011000000110000000000010000",--23276
"000101000000000000000101101011111100",--23277
"111110001000001001010011100000000000",--23278
"001101010110000010110000000000001001",--23279
"001111010110000010000000000000000000",--23280
"111110001110001010000011100000000000",--23281
"111110001100000001110011000000000000",--23282
"111110001010001000110010100000000000",--23283
"001111010110000001110000000000000001",--23284
"111110001010001001110010100000000000",--23285
"111110001100000001010010100000000000",--23286
"111110000110001001000001100000000000",--23287
"001111010110000001000000000000000010",--23288
"111110000110001001000001100000000000",--23289
"111110001010000000110001100000000000",--23290
"011111011011000000110000000000000001",--23291
"111110000110010000010001100000000000",--23292
"001011011000000000110000000000000011",--23293
"101001010100010010100000000000000001",--23294
"010111010101000000000000000010010001",--23295
"001101010100000010110000000101101101",--23296
"001101010110000011000000000000001010",--23297
"001101010110000011010000000000000001",--23298
"001111001110000000110000000000000000",--23299
"001101010110000011100000000000000101",--23300
"001111011100000001000000000000000000",--23301
"111110000110010001000001100000000000",--23302
"001011011000000000110000000000000000",--23303
"001111001110000000110000000000000001",--23304
"001111011100000001000000000000000001",--23305
"111110000110010001000001100000000000",--23306
"001011011000000000110000000000000001",--23307
"001111001110000000110000000000000010",--23308
"001111011100000001000000000000000010",--23309
"111110000110010001000001100000000000",--23310
"001011011000000000110000000000000010",--23311
"011111011011000000100000000000001110",--23312
"001101010110000010110000000000000100",--23313
"001111011000000000110000000000000000",--23314
"001111011000000001000000000000000001",--23315
"001111011000000001010000000000000010",--23316
"001111010110000001100000000000000000",--23317
"111110001100001000110001100000000000",--23318
"001111010110000001100000000000000001",--23319
"111110001100001001000010000000000000",--23320
"111110000110000001000001100000000000",--23321
"001111010110000001000000000000000010",--23322
"111110001000001001010010000000000000",--23323
"111110000110000001000001100000000000",--23324
"001011011000000000110000000000000011",--23325
"000101000000000000000101101101000100",--23326
"010111011011000000100000000000100100",--23327
"001111011000000000110000000000000000",--23328
"001111011000000001000000000000000001",--23329
"001111011000000001010000000000000010",--23330
"111110000110001000110011000000000000",--23331
"001101010110000011100000000000000100",--23332
"001111011100000001110000000000000000",--23333
"111110001100001001110011000000000000",--23334
"111110001000001001000011100000000000",--23335
"001111011100000010000000000000000001",--23336
"111110001110001010000011100000000000",--23337
"111110001100000001110011000000000000",--23338
"111110001010001001010011100000000000",--23339
"001111011100000010000000000000000010",--23340
"111110001110001010000011100000000000",--23341
"111110001100000001110011000000000000",--23342
"001101010110000011100000000000000011",--23343
"011100011101000000000000000000000011",--23344
"101110001101111000000001100000000000",--23345
"011111011011000000110000000000010000",--23346
"000101000000000000000101101101000010",--23347
"111110001000001001010011100000000000",--23348
"001101010110000010110000000000001001",--23349
"001111010110000010000000000000000000",--23350
"111110001110001010000011100000000000",--23351
"111110001100000001110011000000000000",--23352
"111110001010001000110010100000000000",--23353
"001111010110000001110000000000000001",--23354
"111110001010001001110010100000000000",--23355
"111110001100000001010010100000000000",--23356
"111110000110001001000001100000000000",--23357
"001111010110000001000000000000000010",--23358
"111110000110001001000001100000000000",--23359
"111110001010000000110001100000000000",--23360
"011111011011000000110000000000000001",--23361
"111110000110010000010001100000000000",--23362
"001011011000000000110000000000000011",--23363
"101001010100010010100000000000000001",--23364
"010111010101000000000000000001001011",--23365
"001101010100000010110000000101101101",--23366
"001101010110000011000000000000001010",--23367
"001101010110000011010000000000000001",--23368
"001111001110000000110000000000000000",--23369
"001101010110000011100000000000000101",--23370
"001111011100000001000000000000000000",--23371
"111110000110010001000001100000000000",--23372
"001011011000000000110000000000000000",--23373
"001111001110000000110000000000000001",--23374
"001111011100000001000000000000000001",--23375
"111110000110010001000001100000000000",--23376
"001011011000000000110000000000000001",--23377
"001111001110000000110000000000000010",--23378
"001111011100000001000000000000000010",--23379
"111110000110010001000001100000000000",--23380
"001011011000000000110000000000000010",--23381
"011111011011000000100000000000001110",--23382
"001101010110000010110000000000000100",--23383
"001111011000000000110000000000000000",--23384
"001111011000000001000000000000000001",--23385
"001111011000000001010000000000000010",--23386
"001111010110000001100000000000000000",--23387
"111110001100001000110001100000000000",--23388
"001111010110000001100000000000000001",--23389
"111110001100001001000010000000000000",--23390
"111110000110000001000001100000000000",--23391
"001111010110000001000000000000000010",--23392
"111110001000001001010010000000000000",--23393
"111110000110000001000001100000000000",--23394
"001011011000000000110000000000000011",--23395
"000101000000000000000101101110001010",--23396
"010111011011000000100000000000100100",--23397
"001111011000000000110000000000000000",--23398
"001111011000000001000000000000000001",--23399
"001111011000000001010000000000000010",--23400
"111110000110001000110011000000000000",--23401
"001101010110000011100000000000000100",--23402
"001111011100000001110000000000000000",--23403
"111110001100001001110011000000000000",--23404
"111110001000001001000011100000000000",--23405
"001111011100000010000000000000000001",--23406
"111110001110001010000011100000000000",--23407
"111110001100000001110011000000000000",--23408
"111110001010001001010011100000000000",--23409
"001111011100000010000000000000000010",--23410
"111110001110001010000011100000000000",--23411
"111110001100000001110011000000000000",--23412
"001101010110000011100000000000000011",--23413
"011100011101000000000000000000000011",--23414
"101110001101111000000001100000000000",--23415
"011111011011000000110000000000010000",--23416
"000101000000000000000101101110001000",--23417
"111110001000001001010011100000000000",--23418
"001101010110000010110000000000001001",--23419
"001111010110000010000000000000000000",--23420
"111110001110001010000011100000000000",--23421
"111110001100000001110011000000000000",--23422
"111110001010001000110010100000000000",--23423
"001111010110000001110000000000000001",--23424
"111110001010001001110010100000000000",--23425
"111110001100000001010010100000000000",--23426
"111110000110001001000001100000000000",--23427
"001111010110000001000000000000000010",--23428
"111110000110001001000001100000000000",--23429
"111110001010000000110001100000000000",--23430
"011111011011000000110000000000000001",--23431
"111110000110010000010001100000000000",--23432
"001011011000000000110000000000000011",--23433
"101001010100010000100000000000000001",--23434
"101000001111111000000000100000000000",--23435
"001001111100000111111111111111110111",--23436
"101001111100010111100000000000001010",--23437
"000111000000000000000000011001101110",--23438
"101001111100000111100000000000001010",--23439
"001101111100000111111111111111110111",--23440
"101001000000000001000000000001110110",--23441
"001101111100000000011111111111111000",--23442
"001101111100000000101111111111111011",--23443
"001101111100000000111111111111111010",--23444
"001001111100000111111111111111110111",--23445
"101001111100010111100000000000001010",--23446
"000111000000000000000100000011011010",--23447
"101001111100000111100000000000001010",--23448
"001101111100000111111111111111110111",--23449
"001101111100000000011111111111111001",--23450
"010011000011000000010000000011101100",--23451
"001101000000000000100000000011111111",--23452
"001101111100000000111111111111111010",--23453
"001111000110000000110000000000000000",--23454
"001011000000000000110000000100010010",--23455
"001111000110000000110000000000000001",--23456
"001011000000000000110000000100010011",--23457
"001111000110000000110000000000000010",--23458
"001011000000000000110000000100010100",--23459
"001101000000000001000000000110101010",--23460
"101001001000010001000000000000000001",--23461
"001001111100000000101111111111111000",--23462
"010111001001000000000000000011010111",--23463
"001101001000000001010000000101101101",--23464
"001101001010000001100000000000001010",--23465
"001101001010000001110000000000000001",--23466
"001111000110000000110000000000000000",--23467
"001101001010000010000000000000000101",--23468
"001111010000000001000000000000000000",--23469
"111110000110010001000001100000000000",--23470
"001011001100000000110000000000000000",--23471
"001111000110000000110000000000000001",--23472
"001111010000000001000000000000000001",--23473
"111110000110010001000001100000000000",--23474
"001011001100000000110000000000000001",--23475
"001111000110000000110000000000000010",--23476
"001111010000000001000000000000000010",--23477
"111110000110010001000001100000000000",--23478
"001011001100000000110000000000000010",--23479
"011111001111000000100000000000001110",--23480
"001101001010000001010000000000000100",--23481
"001111001100000000110000000000000000",--23482
"001111001100000001000000000000000001",--23483
"001111001100000001010000000000000010",--23484
"001111001010000001100000000000000000",--23485
"111110001100001000110001100000000000",--23486
"001111001010000001100000000000000001",--23487
"111110001100001001000010000000000000",--23488
"111110000110000001000001100000000000",--23489
"001111001010000001000000000000000010",--23490
"111110001000001001010010000000000000",--23491
"111110000110000001000001100000000000",--23492
"001011001100000000110000000000000011",--23493
"000101000000000000000101101111101100",--23494
"010111001111000000100000000000100100",--23495
"001111001100000000110000000000000000",--23496
"001111001100000001000000000000000001",--23497
"001111001100000001010000000000000010",--23498
"111110000110001000110011000000000000",--23499
"001101001010000010000000000000000100",--23500
"001111010000000001110000000000000000",--23501
"111110001100001001110011000000000000",--23502
"111110001000001001000011100000000000",--23503
"001111010000000010000000000000000001",--23504
"111110001110001010000011100000000000",--23505
"111110001100000001110011000000000000",--23506
"111110001010001001010011100000000000",--23507
"001111010000000010000000000000000010",--23508
"111110001110001010000011100000000000",--23509
"111110001100000001110011000000000000",--23510
"001101001010000010000000000000000011",--23511
"011100010001000000000000000000000011",--23512
"101110001101111000000001100000000000",--23513
"011111001111000000110000000000010000",--23514
"000101000000000000000101101111101010",--23515
"111110001000001001010011100000000000",--23516
"001101001010000001010000000000001001",--23517
"001111001010000010000000000000000000",--23518
"111110001110001010000011100000000000",--23519
"111110001100000001110011000000000000",--23520
"111110001010001000110010100000000000",--23521
"001111001010000001110000000000000001",--23522
"111110001010001001110010100000000000",--23523
"111110001100000001010010100000000000",--23524
"111110000110001001000001100000000000",--23525
"001111001010000001000000000000000010",--23526
"111110000110001001000001100000000000",--23527
"111110001010000000110001100000000000",--23528
"011111001111000000110000000000000001",--23529
"111110000110010000010001100000000000",--23530
"001011001100000000110000000000000011",--23531
"101001001000010001000000000000000001",--23532
"010111001001000000000000000010010001",--23533
"001101001000000001010000000101101101",--23534
"001101001010000001100000000000001010",--23535
"001101001010000001110000000000000001",--23536
"001111000110000000110000000000000000",--23537
"001101001010000010000000000000000101",--23538
"001111010000000001000000000000000000",--23539
"111110000110010001000001100000000000",--23540
"001011001100000000110000000000000000",--23541
"001111000110000000110000000000000001",--23542
"001111010000000001000000000000000001",--23543
"111110000110010001000001100000000000",--23544
"001011001100000000110000000000000001",--23545
"001111000110000000110000000000000010",--23546
"001111010000000001000000000000000010",--23547
"111110000110010001000001100000000000",--23548
"001011001100000000110000000000000010",--23549
"011111001111000000100000000000001110",--23550
"001101001010000001010000000000000100",--23551
"001111001100000000110000000000000000",--23552
"001111001100000001000000000000000001",--23553
"001111001100000001010000000000000010",--23554
"001111001010000001100000000000000000",--23555
"111110001100001000110001100000000000",--23556
"001111001010000001100000000000000001",--23557
"111110001100001001000010000000000000",--23558
"111110000110000001000001100000000000",--23559
"001111001010000001000000000000000010",--23560
"111110001000001001010010000000000000",--23561
"111110000110000001000001100000000000",--23562
"001011001100000000110000000000000011",--23563
"000101000000000000000101110000110010",--23564
"010111001111000000100000000000100100",--23565
"001111001100000000110000000000000000",--23566
"001111001100000001000000000000000001",--23567
"001111001100000001010000000000000010",--23568
"111110000110001000110011000000000000",--23569
"001101001010000010000000000000000100",--23570
"001111010000000001110000000000000000",--23571
"111110001100001001110011000000000000",--23572
"111110001000001001000011100000000000",--23573
"001111010000000010000000000000000001",--23574
"111110001110001010000011100000000000",--23575
"111110001100000001110011000000000000",--23576
"111110001010001001010011100000000000",--23577
"001111010000000010000000000000000010",--23578
"111110001110001010000011100000000000",--23579
"111110001100000001110011000000000000",--23580
"001101001010000010000000000000000011",--23581
"011100010001000000000000000000000011",--23582
"101110001101111000000001100000000000",--23583
"011111001111000000110000000000010000",--23584
"000101000000000000000101110000110000",--23585
"111110001000001001010011100000000000",--23586
"001101001010000001010000000000001001",--23587
"001111001010000010000000000000000000",--23588
"111110001110001010000011100000000000",--23589
"111110001100000001110011000000000000",--23590
"111110001010001000110010100000000000",--23591
"001111001010000001110000000000000001",--23592
"111110001010001001110010100000000000",--23593
"111110001100000001010010100000000000",--23594
"111110000110001001000001100000000000",--23595
"001111001010000001000000000000000010",--23596
"111110000110001001000001100000000000",--23597
"111110001010000000110001100000000000",--23598
"011111001111000000110000000000000001",--23599
"111110000110010000010001100000000000",--23600
"001011001100000000110000000000000011",--23601
"101001001000010001000000000000000001",--23602
"010111001001000000000000000001001011",--23603
"001101001000000001010000000101101101",--23604
"001101001010000001100000000000001010",--23605
"001101001010000001110000000000000001",--23606
"001111000110000000110000000000000000",--23607
"001101001010000010000000000000000101",--23608
"001111010000000001000000000000000000",--23609
"111110000110010001000001100000000000",--23610
"001011001100000000110000000000000000",--23611
"001111000110000000110000000000000001",--23612
"001111010000000001000000000000000001",--23613
"111110000110010001000001100000000000",--23614
"001011001100000000110000000000000001",--23615
"001111000110000000110000000000000010",--23616
"001111010000000001000000000000000010",--23617
"111110000110010001000001100000000000",--23618
"001011001100000000110000000000000010",--23619
"011111001111000000100000000000001110",--23620
"001101001010000001010000000000000100",--23621
"001111001100000000110000000000000000",--23622
"001111001100000001000000000000000001",--23623
"001111001100000001010000000000000010",--23624
"001111001010000001100000000000000000",--23625
"111110001100001000110001100000000000",--23626
"001111001010000001100000000000000001",--23627
"111110001100001001000010000000000000",--23628
"111110000110000001000001100000000000",--23629
"001111001010000001000000000000000010",--23630
"111110001000001001010010000000000000",--23631
"111110000110000001000001100000000000",--23632
"001011001100000000110000000000000011",--23633
"000101000000000000000101110001111000",--23634
"010111001111000000100000000000100100",--23635
"001111001100000000110000000000000000",--23636
"001111001100000001000000000000000001",--23637
"001111001100000001010000000000000010",--23638
"111110000110001000110011000000000000",--23639
"001101001010000010000000000000000100",--23640
"001111010000000001110000000000000000",--23641
"111110001100001001110011000000000000",--23642
"111110001000001001000011100000000000",--23643
"001111010000000010000000000000000001",--23644
"111110001110001010000011100000000000",--23645
"111110001100000001110011000000000000",--23646
"111110001010001001010011100000000000",--23647
"001111010000000010000000000000000010",--23648
"111110001110001010000011100000000000",--23649
"111110001100000001110011000000000000",--23650
"001101001010000010000000000000000011",--23651
"011100010001000000000000000000000011",--23652
"101110001101111000000001100000000000",--23653
"011111001111000000110000000000010000",--23654
"000101000000000000000101110001110110",--23655
"111110001000001001010011100000000000",--23656
"001101001010000001010000000000001001",--23657
"001111001010000010000000000000000000",--23658
"111110001110001010000011100000000000",--23659
"111110001100000001110011000000000000",--23660
"111110001010001000110010100000000000",--23661
"001111001010000001110000000000000001",--23662
"111110001010001001110010100000000000",--23663
"111110001100000001010010100000000000",--23664
"111110000110001001000001100000000000",--23665
"001111001010000001000000000000000010",--23666
"111110000110001001000001100000000000",--23667
"111110001010000000110001100000000000",--23668
"011111001111000000110000000000000001",--23669
"111110000110010000010001100000000000",--23670
"001011001100000000110000000000000011",--23671
"101001001000010000100000000000000001",--23672
"101000000111111000000000100000000000",--23673
"001001111100000111111111111111110111",--23674
"101001111100010111100000000000001010",--23675
"000111000000000000000000011001101110",--23676
"101001111100000111100000000000001010",--23677
"001101111100000111111111111111110111",--23678
"101001000000000001000000000001110110",--23679
"001101111100000000011111111111111000",--23680
"001101111100000000101111111111111011",--23681
"001101111100000000111111111111111010",--23682
"001001111100000111111111111111110111",--23683
"101001111100010111100000000000001010",--23684
"000111000000000000000100000011011010",--23685
"101001111100000111100000000000001010",--23686
"001101111100000111111111111111110111",--23687
"001101111100000000011111111111111001",--23688
"010011000011000000100000000011101100",--23689
"001101000000000000100000000100000000",--23690
"001101111100000000111111111111111010",--23691
"001111000110000000110000000000000000",--23692
"001011000000000000110000000100010010",--23693
"001111000110000000110000000000000001",--23694
"001011000000000000110000000100010011",--23695
"001111000110000000110000000000000010",--23696
"001011000000000000110000000100010100",--23697
"001101000000000001000000000110101010",--23698
"101001001000010001000000000000000001",--23699
"001001111100000000101111111111111000",--23700
"010111001001000000000000000011010111",--23701
"001101001000000001010000000101101101",--23702
"001101001010000001100000000000001010",--23703
"001101001010000001110000000000000001",--23704
"001111000110000000110000000000000000",--23705
"001101001010000010000000000000000101",--23706
"001111010000000001000000000000000000",--23707
"111110000110010001000001100000000000",--23708
"001011001100000000110000000000000000",--23709
"001111000110000000110000000000000001",--23710
"001111010000000001000000000000000001",--23711
"111110000110010001000001100000000000",--23712
"001011001100000000110000000000000001",--23713
"001111000110000000110000000000000010",--23714
"001111010000000001000000000000000010",--23715
"111110000110010001000001100000000000",--23716
"001011001100000000110000000000000010",--23717
"011111001111000000100000000000001110",--23718
"001101001010000001010000000000000100",--23719
"001111001100000000110000000000000000",--23720
"001111001100000001000000000000000001",--23721
"001111001100000001010000000000000010",--23722
"001111001010000001100000000000000000",--23723
"111110001100001000110001100000000000",--23724
"001111001010000001100000000000000001",--23725
"111110001100001001000010000000000000",--23726
"111110000110000001000001100000000000",--23727
"001111001010000001000000000000000010",--23728
"111110001000001001010010000000000000",--23729
"111110000110000001000001100000000000",--23730
"001011001100000000110000000000000011",--23731
"000101000000000000000101110011011010",--23732
"010111001111000000100000000000100100",--23733
"001111001100000000110000000000000000",--23734
"001111001100000001000000000000000001",--23735
"001111001100000001010000000000000010",--23736
"111110000110001000110011000000000000",--23737
"001101001010000010000000000000000100",--23738
"001111010000000001110000000000000000",--23739
"111110001100001001110011000000000000",--23740
"111110001000001001000011100000000000",--23741
"001111010000000010000000000000000001",--23742
"111110001110001010000011100000000000",--23743
"111110001100000001110011000000000000",--23744
"111110001010001001010011100000000000",--23745
"001111010000000010000000000000000010",--23746
"111110001110001010000011100000000000",--23747
"111110001100000001110011000000000000",--23748
"001101001010000010000000000000000011",--23749
"011100010001000000000000000000000011",--23750
"101110001101111000000001100000000000",--23751
"011111001111000000110000000000010000",--23752
"000101000000000000000101110011011000",--23753
"111110001000001001010011100000000000",--23754
"001101001010000001010000000000001001",--23755
"001111001010000010000000000000000000",--23756
"111110001110001010000011100000000000",--23757
"111110001100000001110011000000000000",--23758
"111110001010001000110010100000000000",--23759
"001111001010000001110000000000000001",--23760
"111110001010001001110010100000000000",--23761
"111110001100000001010010100000000000",--23762
"111110000110001001000001100000000000",--23763
"001111001010000001000000000000000010",--23764
"111110000110001001000001100000000000",--23765
"111110001010000000110001100000000000",--23766
"011111001111000000110000000000000001",--23767
"111110000110010000010001100000000000",--23768
"001011001100000000110000000000000011",--23769
"101001001000010001000000000000000001",--23770
"010111001001000000000000000010010001",--23771
"001101001000000001010000000101101101",--23772
"001101001010000001100000000000001010",--23773
"001101001010000001110000000000000001",--23774
"001111000110000000110000000000000000",--23775
"001101001010000010000000000000000101",--23776
"001111010000000001000000000000000000",--23777
"111110000110010001000001100000000000",--23778
"001011001100000000110000000000000000",--23779
"001111000110000000110000000000000001",--23780
"001111010000000001000000000000000001",--23781
"111110000110010001000001100000000000",--23782
"001011001100000000110000000000000001",--23783
"001111000110000000110000000000000010",--23784
"001111010000000001000000000000000010",--23785
"111110000110010001000001100000000000",--23786
"001011001100000000110000000000000010",--23787
"011111001111000000100000000000001110",--23788
"001101001010000001010000000000000100",--23789
"001111001100000000110000000000000000",--23790
"001111001100000001000000000000000001",--23791
"001111001100000001010000000000000010",--23792
"001111001010000001100000000000000000",--23793
"111110001100001000110001100000000000",--23794
"001111001010000001100000000000000001",--23795
"111110001100001001000010000000000000",--23796
"111110000110000001000001100000000000",--23797
"001111001010000001000000000000000010",--23798
"111110001000001001010010000000000000",--23799
"111110000110000001000001100000000000",--23800
"001011001100000000110000000000000011",--23801
"000101000000000000000101110100100000",--23802
"010111001111000000100000000000100100",--23803
"001111001100000000110000000000000000",--23804
"001111001100000001000000000000000001",--23805
"001111001100000001010000000000000010",--23806
"111110000110001000110011000000000000",--23807
"001101001010000010000000000000000100",--23808
"001111010000000001110000000000000000",--23809
"111110001100001001110011000000000000",--23810
"111110001000001001000011100000000000",--23811
"001111010000000010000000000000000001",--23812
"111110001110001010000011100000000000",--23813
"111110001100000001110011000000000000",--23814
"111110001010001001010011100000000000",--23815
"001111010000000010000000000000000010",--23816
"111110001110001010000011100000000000",--23817
"111110001100000001110011000000000000",--23818
"001101001010000010000000000000000011",--23819
"011100010001000000000000000000000011",--23820
"101110001101111000000001100000000000",--23821
"011111001111000000110000000000010000",--23822
"000101000000000000000101110100011110",--23823
"111110001000001001010011100000000000",--23824
"001101001010000001010000000000001001",--23825
"001111001010000010000000000000000000",--23826
"111110001110001010000011100000000000",--23827
"111110001100000001110011000000000000",--23828
"111110001010001000110010100000000000",--23829
"001111001010000001110000000000000001",--23830
"111110001010001001110010100000000000",--23831
"111110001100000001010010100000000000",--23832
"111110000110001001000001100000000000",--23833
"001111001010000001000000000000000010",--23834
"111110000110001001000001100000000000",--23835
"111110001010000000110001100000000000",--23836
"011111001111000000110000000000000001",--23837
"111110000110010000010001100000000000",--23838
"001011001100000000110000000000000011",--23839
"101001001000010001000000000000000001",--23840
"010111001001000000000000000001001011",--23841
"001101001000000001010000000101101101",--23842
"001101001010000001100000000000001010",--23843
"001101001010000001110000000000000001",--23844
"001111000110000000110000000000000000",--23845
"001101001010000010000000000000000101",--23846
"001111010000000001000000000000000000",--23847
"111110000110010001000001100000000000",--23848
"001011001100000000110000000000000000",--23849
"001111000110000000110000000000000001",--23850
"001111010000000001000000000000000001",--23851
"111110000110010001000001100000000000",--23852
"001011001100000000110000000000000001",--23853
"001111000110000000110000000000000010",--23854
"001111010000000001000000000000000010",--23855
"111110000110010001000001100000000000",--23856
"001011001100000000110000000000000010",--23857
"011111001111000000100000000000001110",--23858
"001101001010000001010000000000000100",--23859
"001111001100000000110000000000000000",--23860
"001111001100000001000000000000000001",--23861
"001111001100000001010000000000000010",--23862
"001111001010000001100000000000000000",--23863
"111110001100001000110001100000000000",--23864
"001111001010000001100000000000000001",--23865
"111110001100001001000010000000000000",--23866
"111110000110000001000001100000000000",--23867
"001111001010000001000000000000000010",--23868
"111110001000001001010010000000000000",--23869
"111110000110000001000001100000000000",--23870
"001011001100000000110000000000000011",--23871
"000101000000000000000101110101100110",--23872
"010111001111000000100000000000100100",--23873
"001111001100000000110000000000000000",--23874
"001111001100000001000000000000000001",--23875
"001111001100000001010000000000000010",--23876
"111110000110001000110011000000000000",--23877
"001101001010000010000000000000000100",--23878
"001111010000000001110000000000000000",--23879
"111110001100001001110011000000000000",--23880
"111110001000001001000011100000000000",--23881
"001111010000000010000000000000000001",--23882
"111110001110001010000011100000000000",--23883
"111110001100000001110011000000000000",--23884
"111110001010001001010011100000000000",--23885
"001111010000000010000000000000000010",--23886
"111110001110001010000011100000000000",--23887
"111110001100000001110011000000000000",--23888
"001101001010000010000000000000000011",--23889
"011100010001000000000000000000000011",--23890
"101110001101111000000001100000000000",--23891
"011111001111000000110000000000010000",--23892
"000101000000000000000101110101100100",--23893
"111110001000001001010011100000000000",--23894
"001101001010000001010000000000001001",--23895
"001111001010000010000000000000000000",--23896
"111110001110001010000011100000000000",--23897
"111110001100000001110011000000000000",--23898
"111110001010001000110010100000000000",--23899
"001111001010000001110000000000000001",--23900
"111110001010001001110010100000000000",--23901
"111110001100000001010010100000000000",--23902
"111110000110001001000001100000000000",--23903
"001111001010000001000000000000000010",--23904
"111110000110001001000001100000000000",--23905
"111110001010000000110001100000000000",--23906
"011111001111000000110000000000000001",--23907
"111110000110010000010001100000000000",--23908
"001011001100000000110000000000000011",--23909
"101001001000010000100000000000000001",--23910
"101000000111111000000000100000000000",--23911
"001001111100000111111111111111110111",--23912
"101001111100010111100000000000001010",--23913
"000111000000000000000000011001101110",--23914
"101001111100000111100000000000001010",--23915
"001101111100000111111111111111110111",--23916
"101001000000000001000000000001110110",--23917
"001101111100000000011111111111111000",--23918
"001101111100000000101111111111111011",--23919
"001101111100000000111111111111111010",--23920
"001001111100000111111111111111110111",--23921
"101001111100010111100000000000001010",--23922
"000111000000000000000100000011011010",--23923
"101001111100000111100000000000001010",--23924
"001101111100000111111111111111110111",--23925
"001101111100000000011111111111111001",--23926
"010011000011000000110000000011101100",--23927
"001101000000000000100000000100000001",--23928
"001101111100000000111111111111111010",--23929
"001111000110000000110000000000000000",--23930
"001011000000000000110000000100010010",--23931
"001111000110000000110000000000000001",--23932
"001011000000000000110000000100010011",--23933
"001111000110000000110000000000000010",--23934
"001011000000000000110000000100010100",--23935
"001101000000000001000000000110101010",--23936
"101001001000010001000000000000000001",--23937
"001001111100000000101111111111111000",--23938
"010111001001000000000000000011010111",--23939
"001101001000000001010000000101101101",--23940
"001101001010000001100000000000001010",--23941
"001101001010000001110000000000000001",--23942
"001111000110000000110000000000000000",--23943
"001101001010000010000000000000000101",--23944
"001111010000000001000000000000000000",--23945
"111110000110010001000001100000000000",--23946
"001011001100000000110000000000000000",--23947
"001111000110000000110000000000000001",--23948
"001111010000000001000000000000000001",--23949
"111110000110010001000001100000000000",--23950
"001011001100000000110000000000000001",--23951
"001111000110000000110000000000000010",--23952
"001111010000000001000000000000000010",--23953
"111110000110010001000001100000000000",--23954
"001011001100000000110000000000000010",--23955
"011111001111000000100000000000001110",--23956
"001101001010000001010000000000000100",--23957
"001111001100000000110000000000000000",--23958
"001111001100000001000000000000000001",--23959
"001111001100000001010000000000000010",--23960
"001111001010000001100000000000000000",--23961
"111110001100001000110001100000000000",--23962
"001111001010000001100000000000000001",--23963
"111110001100001001000010000000000000",--23964
"111110000110000001000001100000000000",--23965
"001111001010000001000000000000000010",--23966
"111110001000001001010010000000000000",--23967
"111110000110000001000001100000000000",--23968
"001011001100000000110000000000000011",--23969
"000101000000000000000101110111001000",--23970
"010111001111000000100000000000100100",--23971
"001111001100000000110000000000000000",--23972
"001111001100000001000000000000000001",--23973
"001111001100000001010000000000000010",--23974
"111110000110001000110011000000000000",--23975
"001101001010000010000000000000000100",--23976
"001111010000000001110000000000000000",--23977
"111110001100001001110011000000000000",--23978
"111110001000001001000011100000000000",--23979
"001111010000000010000000000000000001",--23980
"111110001110001010000011100000000000",--23981
"111110001100000001110011000000000000",--23982
"111110001010001001010011100000000000",--23983
"001111010000000010000000000000000010",--23984
"111110001110001010000011100000000000",--23985
"111110001100000001110011000000000000",--23986
"001101001010000010000000000000000011",--23987
"011100010001000000000000000000000011",--23988
"101110001101111000000001100000000000",--23989
"011111001111000000110000000000010000",--23990
"000101000000000000000101110111000110",--23991
"111110001000001001010011100000000000",--23992
"001101001010000001010000000000001001",--23993
"001111001010000010000000000000000000",--23994
"111110001110001010000011100000000000",--23995
"111110001100000001110011000000000000",--23996
"111110001010001000110010100000000000",--23997
"001111001010000001110000000000000001",--23998
"111110001010001001110010100000000000",--23999
"111110001100000001010010100000000000",--24000
"111110000110001001000001100000000000",--24001
"001111001010000001000000000000000010",--24002
"111110000110001001000001100000000000",--24003
"111110001010000000110001100000000000",--24004
"011111001111000000110000000000000001",--24005
"111110000110010000010001100000000000",--24006
"001011001100000000110000000000000011",--24007
"101001001000010001000000000000000001",--24008
"010111001001000000000000000010010001",--24009
"001101001000000001010000000101101101",--24010
"001101001010000001100000000000001010",--24011
"001101001010000001110000000000000001",--24012
"001111000110000000110000000000000000",--24013
"001101001010000010000000000000000101",--24014
"001111010000000001000000000000000000",--24015
"111110000110010001000001100000000000",--24016
"001011001100000000110000000000000000",--24017
"001111000110000000110000000000000001",--24018
"001111010000000001000000000000000001",--24019
"111110000110010001000001100000000000",--24020
"001011001100000000110000000000000001",--24021
"001111000110000000110000000000000010",--24022
"001111010000000001000000000000000010",--24023
"111110000110010001000001100000000000",--24024
"001011001100000000110000000000000010",--24025
"011111001111000000100000000000001110",--24026
"001101001010000001010000000000000100",--24027
"001111001100000000110000000000000000",--24028
"001111001100000001000000000000000001",--24029
"001111001100000001010000000000000010",--24030
"001111001010000001100000000000000000",--24031
"111110001100001000110001100000000000",--24032
"001111001010000001100000000000000001",--24033
"111110001100001001000010000000000000",--24034
"111110000110000001000001100000000000",--24035
"001111001010000001000000000000000010",--24036
"111110001000001001010010000000000000",--24037
"111110000110000001000001100000000000",--24038
"001011001100000000110000000000000011",--24039
"000101000000000000000101111000001110",--24040
"010111001111000000100000000000100100",--24041
"001111001100000000110000000000000000",--24042
"001111001100000001000000000000000001",--24043
"001111001100000001010000000000000010",--24044
"111110000110001000110011000000000000",--24045
"001101001010000010000000000000000100",--24046
"001111010000000001110000000000000000",--24047
"111110001100001001110011000000000000",--24048
"111110001000001001000011100000000000",--24049
"001111010000000010000000000000000001",--24050
"111110001110001010000011100000000000",--24051
"111110001100000001110011000000000000",--24052
"111110001010001001010011100000000000",--24053
"001111010000000010000000000000000010",--24054
"111110001110001010000011100000000000",--24055
"111110001100000001110011000000000000",--24056
"001101001010000010000000000000000011",--24057
"011100010001000000000000000000000011",--24058
"101110001101111000000001100000000000",--24059
"011111001111000000110000000000010000",--24060
"000101000000000000000101111000001100",--24061
"111110001000001001010011100000000000",--24062
"001101001010000001010000000000001001",--24063
"001111001010000010000000000000000000",--24064
"111110001110001010000011100000000000",--24065
"111110001100000001110011000000000000",--24066
"111110001010001000110010100000000000",--24067
"001111001010000001110000000000000001",--24068
"111110001010001001110010100000000000",--24069
"111110001100000001010010100000000000",--24070
"111110000110001001000001100000000000",--24071
"001111001010000001000000000000000010",--24072
"111110000110001001000001100000000000",--24073
"111110001010000000110001100000000000",--24074
"011111001111000000110000000000000001",--24075
"111110000110010000010001100000000000",--24076
"001011001100000000110000000000000011",--24077
"101001001000010001000000000000000001",--24078
"010111001001000000000000000001001011",--24079
"001101001000000001010000000101101101",--24080
"001101001010000001100000000000001010",--24081
"001101001010000001110000000000000001",--24082
"001111000110000000110000000000000000",--24083
"001101001010000010000000000000000101",--24084
"001111010000000001000000000000000000",--24085
"111110000110010001000001100000000000",--24086
"001011001100000000110000000000000000",--24087
"001111000110000000110000000000000001",--24088
"001111010000000001000000000000000001",--24089
"111110000110010001000001100000000000",--24090
"001011001100000000110000000000000001",--24091
"001111000110000000110000000000000010",--24092
"001111010000000001000000000000000010",--24093
"111110000110010001000001100000000000",--24094
"001011001100000000110000000000000010",--24095
"011111001111000000100000000000001110",--24096
"001101001010000001010000000000000100",--24097
"001111001100000000110000000000000000",--24098
"001111001100000001000000000000000001",--24099
"001111001100000001010000000000000010",--24100
"001111001010000001100000000000000000",--24101
"111110001100001000110001100000000000",--24102
"001111001010000001100000000000000001",--24103
"111110001100001001000010000000000000",--24104
"111110000110000001000001100000000000",--24105
"001111001010000001000000000000000010",--24106
"111110001000001001010010000000000000",--24107
"111110000110000001000001100000000000",--24108
"001011001100000000110000000000000011",--24109
"000101000000000000000101111001010100",--24110
"010111001111000000100000000000100100",--24111
"001111001100000000110000000000000000",--24112
"001111001100000001000000000000000001",--24113
"001111001100000001010000000000000010",--24114
"111110000110001000110011000000000000",--24115
"001101001010000010000000000000000100",--24116
"001111010000000001110000000000000000",--24117
"111110001100001001110011000000000000",--24118
"111110001000001001000011100000000000",--24119
"001111010000000010000000000000000001",--24120
"111110001110001010000011100000000000",--24121
"111110001100000001110011000000000000",--24122
"111110001010001001010011100000000000",--24123
"001111010000000010000000000000000010",--24124
"111110001110001010000011100000000000",--24125
"111110001100000001110011000000000000",--24126
"001101001010000010000000000000000011",--24127
"011100010001000000000000000000000011",--24128
"101110001101111000000001100000000000",--24129
"011111001111000000110000000000010000",--24130
"000101000000000000000101111001010010",--24131
"111110001000001001010011100000000000",--24132
"001101001010000001010000000000001001",--24133
"001111001010000010000000000000000000",--24134
"111110001110001010000011100000000000",--24135
"111110001100000001110011000000000000",--24136
"111110001010001000110010100000000000",--24137
"001111001010000001110000000000000001",--24138
"111110001010001001110010100000000000",--24139
"111110001100000001010010100000000000",--24140
"111110000110001001000001100000000000",--24141
"001111001010000001000000000000000010",--24142
"111110000110001001000001100000000000",--24143
"111110001010000000110001100000000000",--24144
"011111001111000000110000000000000001",--24145
"111110000110010000010001100000000000",--24146
"001011001100000000110000000000000011",--24147
"101001001000010000100000000000000001",--24148
"101000000111111000000000100000000000",--24149
"001001111100000111111111111111110111",--24150
"101001111100010111100000000000001010",--24151
"000111000000000000000000011001101110",--24152
"101001111100000111100000000000001010",--24153
"001101111100000111111111111111110111",--24154
"101001000000000001000000000001110110",--24155
"001101111100000000011111111111111000",--24156
"001101111100000000101111111111111011",--24157
"001101111100000000111111111111111010",--24158
"001001111100000111111111111111110111",--24159
"101001111100010111100000000000001010",--24160
"000111000000000000000100000011011010",--24161
"101001111100000111100000000000001010",--24162
"001101111100000111111111111111110111",--24163
"001101111100000000011111111111111001",--24164
"010011000011000001000000000011101100",--24165
"001101000000000000010000000100000010",--24166
"001101111100000000111111111111111010",--24167
"001111000110000000110000000000000000",--24168
"001011000000000000110000000100010010",--24169
"001111000110000000110000000000000001",--24170
"001011000000000000110000000100010011",--24171
"001111000110000000110000000000000010",--24172
"001011000000000000110000000100010100",--24173
"001101000000000000100000000110101010",--24174
"101001000100010000100000000000000001",--24175
"001001111100000000011111111111111000",--24176
"010111000101000000000000000011010111",--24177
"001101000100000001000000000101101101",--24178
"001101001000000001010000000000001010",--24179
"001101001000000001100000000000000001",--24180
"001111000110000000110000000000000000",--24181
"001101001000000001110000000000000101",--24182
"001111001110000001000000000000000000",--24183
"111110000110010001000001100000000000",--24184
"001011001010000000110000000000000000",--24185
"001111000110000000110000000000000001",--24186
"001111001110000001000000000000000001",--24187
"111110000110010001000001100000000000",--24188
"001011001010000000110000000000000001",--24189
"001111000110000000110000000000000010",--24190
"001111001110000001000000000000000010",--24191
"111110000110010001000001100000000000",--24192
"001011001010000000110000000000000010",--24193
"011111001101000000100000000000001110",--24194
"001101001000000001000000000000000100",--24195
"001111001010000000110000000000000000",--24196
"001111001010000001000000000000000001",--24197
"001111001010000001010000000000000010",--24198
"001111001000000001100000000000000000",--24199
"111110001100001000110001100000000000",--24200
"001111001000000001100000000000000001",--24201
"111110001100001001000010000000000000",--24202
"111110000110000001000001100000000000",--24203
"001111001000000001000000000000000010",--24204
"111110001000001001010010000000000000",--24205
"111110000110000001000001100000000000",--24206
"001011001010000000110000000000000011",--24207
"000101000000000000000101111010110110",--24208
"010111001101000000100000000000100100",--24209
"001111001010000000110000000000000000",--24210
"001111001010000001000000000000000001",--24211
"001111001010000001010000000000000010",--24212
"111110000110001000110011000000000000",--24213
"001101001000000001110000000000000100",--24214
"001111001110000001110000000000000000",--24215
"111110001100001001110011000000000000",--24216
"111110001000001001000011100000000000",--24217
"001111001110000010000000000000000001",--24218
"111110001110001010000011100000000000",--24219
"111110001100000001110011000000000000",--24220
"111110001010001001010011100000000000",--24221
"001111001110000010000000000000000010",--24222
"111110001110001010000011100000000000",--24223
"111110001100000001110011000000000000",--24224
"001101001000000001110000000000000011",--24225
"011100001111000000000000000000000011",--24226
"101110001101111000000001100000000000",--24227
"011111001101000000110000000000010000",--24228
"000101000000000000000101111010110100",--24229
"111110001000001001010011100000000000",--24230
"001101001000000001000000000000001001",--24231
"001111001000000010000000000000000000",--24232
"111110001110001010000011100000000000",--24233
"111110001100000001110011000000000000",--24234
"111110001010001000110010100000000000",--24235
"001111001000000001110000000000000001",--24236
"111110001010001001110010100000000000",--24237
"111110001100000001010010100000000000",--24238
"111110000110001001000001100000000000",--24239
"001111001000000001000000000000000010",--24240
"111110000110001001000001100000000000",--24241
"111110001010000000110001100000000000",--24242
"011111001101000000110000000000000001",--24243
"111110000110010000010001100000000000",--24244
"001011001010000000110000000000000011",--24245
"101001000100010000100000000000000001",--24246
"010111000101000000000000000010010001",--24247
"001101000100000001000000000101101101",--24248
"001101001000000001010000000000001010",--24249
"001101001000000001100000000000000001",--24250
"001111000110000000110000000000000000",--24251
"001101001000000001110000000000000101",--24252
"001111001110000001000000000000000000",--24253
"111110000110010001000001100000000000",--24254
"001011001010000000110000000000000000",--24255
"001111000110000000110000000000000001",--24256
"001111001110000001000000000000000001",--24257
"111110000110010001000001100000000000",--24258
"001011001010000000110000000000000001",--24259
"001111000110000000110000000000000010",--24260
"001111001110000001000000000000000010",--24261
"111110000110010001000001100000000000",--24262
"001011001010000000110000000000000010",--24263
"011111001101000000100000000000001110",--24264
"001101001000000001000000000000000100",--24265
"001111001010000000110000000000000000",--24266
"001111001010000001000000000000000001",--24267
"001111001010000001010000000000000010",--24268
"001111001000000001100000000000000000",--24269
"111110001100001000110001100000000000",--24270
"001111001000000001100000000000000001",--24271
"111110001100001001000010000000000000",--24272
"111110000110000001000001100000000000",--24273
"001111001000000001000000000000000010",--24274
"111110001000001001010010000000000000",--24275
"111110000110000001000001100000000000",--24276
"001011001010000000110000000000000011",--24277
"000101000000000000000101111011111100",--24278
"010111001101000000100000000000100100",--24279
"001111001010000000110000000000000000",--24280
"001111001010000001000000000000000001",--24281
"001111001010000001010000000000000010",--24282
"111110000110001000110011000000000000",--24283
"001101001000000001110000000000000100",--24284
"001111001110000001110000000000000000",--24285
"111110001100001001110011000000000000",--24286
"111110001000001001000011100000000000",--24287
"001111001110000010000000000000000001",--24288
"111110001110001010000011100000000000",--24289
"111110001100000001110011000000000000",--24290
"111110001010001001010011100000000000",--24291
"001111001110000010000000000000000010",--24292
"111110001110001010000011100000000000",--24293
"111110001100000001110011000000000000",--24294
"001101001000000001110000000000000011",--24295
"011100001111000000000000000000000011",--24296
"101110001101111000000001100000000000",--24297
"011111001101000000110000000000010000",--24298
"000101000000000000000101111011111010",--24299
"111110001000001001010011100000000000",--24300
"001101001000000001000000000000001001",--24301
"001111001000000010000000000000000000",--24302
"111110001110001010000011100000000000",--24303
"111110001100000001110011000000000000",--24304
"111110001010001000110010100000000000",--24305
"001111001000000001110000000000000001",--24306
"111110001010001001110010100000000000",--24307
"111110001100000001010010100000000000",--24308
"111110000110001001000001100000000000",--24309
"001111001000000001000000000000000010",--24310
"111110000110001001000001100000000000",--24311
"111110001010000000110001100000000000",--24312
"011111001101000000110000000000000001",--24313
"111110000110010000010001100000000000",--24314
"001011001010000000110000000000000011",--24315
"101001000100010000100000000000000001",--24316
"010111000101000000000000000001001011",--24317
"001101000100000001000000000101101101",--24318
"001101001000000001010000000000001010",--24319
"001101001000000001100000000000000001",--24320
"001111000110000000110000000000000000",--24321
"001101001000000001110000000000000101",--24322
"001111001110000001000000000000000000",--24323
"111110000110010001000001100000000000",--24324
"001011001010000000110000000000000000",--24325
"001111000110000000110000000000000001",--24326
"001111001110000001000000000000000001",--24327
"111110000110010001000001100000000000",--24328
"001011001010000000110000000000000001",--24329
"001111000110000000110000000000000010",--24330
"001111001110000001000000000000000010",--24331
"111110000110010001000001100000000000",--24332
"001011001010000000110000000000000010",--24333
"011111001101000000100000000000001110",--24334
"001101001000000001000000000000000100",--24335
"001111001010000000110000000000000000",--24336
"001111001010000001000000000000000001",--24337
"001111001010000001010000000000000010",--24338
"001111001000000001100000000000000000",--24339
"111110001100001000110001100000000000",--24340
"001111001000000001100000000000000001",--24341
"111110001100001001000010000000000000",--24342
"111110000110000001000001100000000000",--24343
"001111001000000001000000000000000010",--24344
"111110001000001001010010000000000000",--24345
"111110000110000001000001100000000000",--24346
"001011001010000000110000000000000011",--24347
"000101000000000000000101111101000010",--24348
"010111001101000000100000000000100100",--24349
"001111001010000000110000000000000000",--24350
"001111001010000001000000000000000001",--24351
"001111001010000001010000000000000010",--24352
"111110000110001000110011000000000000",--24353
"001101001000000001110000000000000100",--24354
"001111001110000001110000000000000000",--24355
"111110001100001001110011000000000000",--24356
"111110001000001001000011100000000000",--24357
"001111001110000010000000000000000001",--24358
"111110001110001010000011100000000000",--24359
"111110001100000001110011000000000000",--24360
"111110001010001001010011100000000000",--24361
"001111001110000010000000000000000010",--24362
"111110001110001010000011100000000000",--24363
"111110001100000001110011000000000000",--24364
"001101001000000001110000000000000011",--24365
"011100001111000000000000000000000011",--24366
"101110001101111000000001100000000000",--24367
"011111001101000000110000000000010000",--24368
"000101000000000000000101111101000000",--24369
"111110001000001001010011100000000000",--24370
"001101001000000001000000000000001001",--24371
"001111001000000010000000000000000000",--24372
"111110001110001010000011100000000000",--24373
"111110001100000001110011000000000000",--24374
"111110001010001000110010100000000000",--24375
"001111001000000001110000000000000001",--24376
"111110001010001001110010100000000000",--24377
"111110001100000001010010100000000000",--24378
"111110000110001001000001100000000000",--24379
"001111001000000001000000000000000010",--24380
"111110000110001001000001100000000000",--24381
"111110001010000000110001100000000000",--24382
"011111001101000000110000000000000001",--24383
"111110000110010000010001100000000000",--24384
"001011001010000000110000000000000011",--24385
"101001000100010000100000000000000001",--24386
"101000000111111000000000100000000000",--24387
"001001111100000111111111111111110111",--24388
"101001111100010111100000000000001010",--24389
"000111000000000000000000011001101110",--24390
"101001111100000111100000000000001010",--24391
"001101111100000111111111111111110111",--24392
"101001000000000001000000000001110110",--24393
"001101111100000000011111111111111000",--24394
"001101111100000000101111111111111011",--24395
"001101111100000000111111111111111010",--24396
"001001111100000111111111111111110111",--24397
"101001111100010111100000000000001010",--24398
"000111000000000000000100000011011010",--24399
"101001111100000111100000000000001010",--24400
"001101111100000111111111111111110111",--24401
"001101111100000000011111111111111101",--24402
"001101111100000000111111111111111100",--24403
"001100000110000000010001000000000000",--24404
"001111000000000000110000000100011101",--24405
"001111000100000001000000000000000000",--24406
"001111000000000001010000000100100000",--24407
"111110001000001001010010000000000000",--24408
"111110000110000001000001100000000000",--24409
"001011000000000000110000000100011101",--24410
"001111000000000000110000000100011110",--24411
"001111000100000001000000000000000001",--24412
"001111000000000001010000000100100001",--24413
"111110001000001001010010000000000000",--24414
"111110000110000001000001100000000000",--24415
"001011000000000000110000000100011110",--24416
"001111000000000000110000000100011111",--24417
"001111000100000001000000000000000010",--24418
"001111000000000001010000000100100010",--24419
"111110001000001001010010000000000000",--24420
"111110000110000001000001100000000000",--24421
"001011000000000000110000000100011111",--24422
"001101111100000000011111111111111101",--24423
"101001000010000000010000000000000001",--24424
"011011000010000001011111100000000000",--24425
"001101111100000000111111111111111110",--24426
"001100000110000000010001000000000000",--24427
"010111000100000000001111100000000000",--24428
"001101111100000001001111111111111111",--24429
"001100001000000000010001000000000000",--24430
"010000000101000000000000000001011011",--24431
"001101111100000000100000000000000000",--24432
"001101000100000001010000000000000101",--24433
"001101000100000001100000000000000111",--24434
"001101000100000001110000000000000001",--24435
"001101000100000010000000000000000100",--24436
"001100001010000000010010100000000000",--24437
"001111001010000000110000000000000000",--24438
"001011000000000000110000000100100000",--24439
"001111001010000000110000000000000001",--24440
"001011000000000000110000000100100001",--24441
"001111001010000000110000000000000010",--24442
"001011000000000000110000000100100010",--24443
"001101000100000001010000000000000110",--24444
"001101001010000001010000000000000000",--24445
"001100001100000000010011000000000000",--24446
"001100001110000000010011100000000000",--24447
"001001111100000010001111111111111100",--24448
"001001111100000000011111111111111011",--24449
"001001111100000001111111111111111010",--24450
"001001111100000001101111111111111001",--24451
"001001111100000001011111111111111000",--24452
"010000001011000000000000000000001000",--24453
"001101000000000000010000000011111110",--24454
"101000001111111000000001100000000000",--24455
"101000001101111000000001000000000000",--24456
"001001111100000111111111111111110111",--24457
"101001111100010111100000000000001010",--24458
"000111000000000000000100101110010000",--24459
"101001111100000111100000000000001010",--24460
"001101111100000111111111111111110111",--24461
"001101111100000000011111111111111000",--24462
"010011000011000000010000000000001000",--24463
"001101000000000000010000000011111111",--24464
"001101111100000000101111111111111001",--24465
"001101111100000000111111111111111010",--24466
"001001111100000111111111111111110111",--24467
"101001111100010111100000000000001010",--24468
"000111000000000000000100101110010000",--24469
"101001111100000111100000000000001010",--24470
"001101111100000111111111111111110111",--24471
"001101111100000000011111111111111000",--24472
"010011000011000000100000000000001000",--24473
"001101000000000000010000000100000000",--24474
"001101111100000000101111111111111001",--24475
"001101111100000000111111111111111010",--24476
"001001111100000111111111111111110111",--24477
"101001111100010111100000000000001010",--24478
"000111000000000000000100101110010000",--24479
"101001111100000111100000000000001010",--24480
"001101111100000111111111111111110111",--24481
"001101111100000000011111111111111000",--24482
"010011000011000000110000000000001000",--24483
"001101000000000000010000000100000001",--24484
"001101111100000000101111111111111001",--24485
"001101111100000000111111111111111010",--24486
"001001111100000111111111111111110111",--24487
"101001111100010111100000000000001010",--24488
"000111000000000000000100101110010000",--24489
"101001111100000111100000000000001010",--24490
"001101111100000111111111111111110111",--24491
"001101111100000000011111111111111000",--24492
"010011000011000001000000000000001000",--24493
"001101000000000000010000000100000010",--24494
"001101111100000000101111111111111001",--24495
"001101111100000000111111111111111010",--24496
"001001111100000111111111111111110111",--24497
"101001111100010111100000000000001010",--24498
"000111000000000000000100101110010000",--24499
"101001111100000111100000000000001010",--24500
"001101111100000111111111111111110111",--24501
"001101111100000000011111111111111011",--24502
"001101111100000000111111111111111100",--24503
"001100000110000000010001000000000000",--24504
"001111000000000000110000000100011101",--24505
"001111000100000001000000000000000000",--24506
"001111000000000001010000000100100000",--24507
"111110001000001001010010000000000000",--24508
"111110000110000001000001100000000000",--24509
"001011000000000000110000000100011101",--24510
"001111000000000000110000000100011110",--24511
"001111000100000001000000000000000001",--24512
"001111000000000001010000000100100001",--24513
"111110001000001001010010000000000000",--24514
"111110000110000001000001100000000000",--24515
"001011000000000000110000000100011110",--24516
"001111000000000000110000000100011111",--24517
"001111000100000001000000000000000010",--24518
"001111000000000001010000000100100010",--24519
"111110001000001001010010000000000000",--24520
"111110000110000001000001100000000000",--24521
"001011000000000000110000000100011111",--24522
"101001000010000000010000000000000001",--24523
"011011000010000001011111100000000000",--24524
"001101111100000000111111111111111110",--24525
"001100000110000000010001000000000000",--24526
"010111000100000000001111100000000000",--24527
"001101111100000001001111111111111111",--24528
"001100001000000000010001000000000000",--24529
"010000000101000000000000000000101101",--24530
"001101111100000000100000000000000000",--24531
"001101000100000001010000000000000101",--24532
"001101000100000001100000000000000111",--24533
"001101000100000001110000000000000001",--24534
"001101000100000010000000000000000100",--24535
"001100001010000000010010100000000000",--24536
"001111001010000000110000000000000000",--24537
"001011000000000000110000000100100000",--24538
"001111001010000000110000000000000001",--24539
"001011000000000000110000000100100001",--24540
"001111001010000000110000000000000010",--24541
"001011000000000000110000000100100010",--24542
"001101000100000001010000000000000110",--24543
"001101001010000001010000000000000000",--24544
"001100001100000000010001000000000000",--24545
"001100001110000000010001100000000000",--24546
"001001111100000010001111111111111100",--24547
"001001111100000000011111111111111011",--24548
"101000001011111000000000100000000000",--24549
"001001111100000111111111111111111010",--24550
"101001111100010111100000000000000111",--24551
"000111000000000000000101000111001101",--24552
"101001111100000111100000000000000111",--24553
"001101111100000111111111111111111010",--24554
"001101111100000000011111111111111011",--24555
"001101111100000000111111111111111100",--24556
"001100000110000000010001000000000000",--24557
"001111000000000000110000000100011101",--24558
"001111000100000001000000000000000000",--24559
"001111000000000001010000000100100000",--24560
"111110001000001001010010000000000000",--24561
"111110000110000001000001100000000000",--24562
"001011000000000000110000000100011101",--24563
"001111000000000000110000000100011110",--24564
"001111000100000001000000000000000001",--24565
"001111000000000001010000000100100001",--24566
"111110001000001001010010000000000000",--24567
"111110000110000001000001100000000000",--24568
"001011000000000000110000000100011110",--24569
"001111000000000000110000000100011111",--24570
"001111000100000001000000000000000010",--24571
"001111000000000001010000000100100010",--24572
"111110001000001001010010000000000000",--24573
"111110000110000001000001100000000000",--24574
"001011000000000000110000000100011111",--24575
"101001000010000000100000000000000001",--24576
"011011000100000001011111100000000000",--24577
"001101111100000000111111111111111110",--24578
"001100000110000000100000100000000000",--24579
"010111000010000000001111100000000000",--24580
"001101111100000000111111111111111111",--24581
"001100000110000000100000100000000000",--24582
"001001111100000000101111111111111100",--24583
"010000000011000000000000000000000110",--24584
"001101111100000000010000000000000000",--24585
"001001111100000111111111111111111011",--24586
"101001111100010111100000000000000110",--24587
"000111000000000000000101011001110000",--24588
"101001111100000111100000000000000110",--24589
"001101111100000111111111111111111011",--24590
"001101111100000000011111111111111100",--24591
"101001000010000000100000000000000001",--24592
"001101111100000000010000000000000000",--24593
"011011000100000001011111100000000000",--24594
"000101000000000000000101101010010001",--24595
"011011001100000001011111100000000000",--24596
"001100001000000000010011100000000000",--24597
"001101001110000010000000000000000010",--24598
"001100010000000001100100000000000000",--24599
"010111010000000000001111100000000000",--24600
"001100001000000000010100000000000000",--24601
"001101010000000010000000000000000010",--24602
"001100010000000001100100000000000000",--24603
"001100000110000000010100100000000000",--24604
"001101010010000010010000000000000010",--24605
"001100010010000001100100100000000000",--24606
"011100010011000010000000000000010100",--24607
"001100001010000000010100100000000000",--24608
"001101010010000010010000000000000010",--24609
"001100010010000001100100100000000000",--24610
"011100010011000010000000000000001110",--24611
"101001000010010010010000000000000001",--24612
"001100001000000010010100100000000000",--24613
"001101010010000010010000000000000010",--24614
"001100010010000001100100100000000000",--24615
"011100010011000010000000000000000111",--24616
"101001000010000010010000000000000001",--24617
"001100001000000010010100100000000000",--24618
"001101010010000010010000000000000010",--24619
"001100010010000001100100100000000000",--24620
"010000010011000010000000000010110101",--24621
"011011001100000001011111100000000000",--24622
"000101000000000000000110000000110101",--24623
"011011001100000001011111100000000000",--24624
"000101000000000000000110000000110101",--24625
"011011001100000001011111100000000000",--24626
"000101000000000000000110000000110101",--24627
"011011001100000001011111100000000000",--24628
"001100001000000000010000100000000000",--24629
"001101000010000000100000000000000010",--24630
"001100000100000001100001100000000000",--24631
"010111000110000000001111100000000000",--24632
"001101000010000000110000000000000011",--24633
"001100000110000001100010000000000000",--24634
"001001111100000000010000000000000000",--24635
"001001111100000000111111111111111111",--24636
"001001111100000000101111111111111110",--24637
"001001111100000001101111111111111101",--24638
"010000001001000000000000000001011001",--24639
"001101000010000001000000000000000101",--24640
"001101000010000001010000000000000111",--24641
"001101000010000001110000000000000001",--24642
"001101000010000010000000000000000100",--24643
"001100001000000001100010000000000000",--24644
"001111001000000000110000000000000000",--24645
"001011000000000000110000000100100000",--24646
"001111001000000000110000000000000001",--24647
"001011000000000000110000000100100001",--24648
"001111001000000000110000000000000010",--24649
"001011000000000000110000000100100010",--24650
"001101000010000001000000000000000110",--24651
"001101001000000001000000000000000000",--24652
"001100001010000001100010100000000000",--24653
"001100001110000001100011100000000000",--24654
"001001111100000010001111111111111100",--24655
"001001111100000001111111111111111011",--24656
"001001111100000001011111111111111010",--24657
"001001111100000001001111111111111001",--24658
"010000001001000000000000000000001000",--24659
"001101000000000000010000000011111110",--24660
"101000001111111000000001100000000000",--24661
"101000001011111000000001000000000000",--24662
"001001111100000111111111111111111000",--24663
"101001111100010111100000000000001001",--24664
"000111000000000000000100101110010000",--24665
"101001111100000111100000000000001001",--24666
"001101111100000111111111111111111000",--24667
"001101111100000000011111111111111001",--24668
"010011000011000000010000000000001000",--24669
"001101000000000000010000000011111111",--24670
"001101111100000000101111111111111010",--24671
"001101111100000000111111111111111011",--24672
"001001111100000111111111111111111000",--24673
"101001111100010111100000000000001001",--24674
"000111000000000000000100101110010000",--24675
"101001111100000111100000000000001001",--24676
"001101111100000111111111111111111000",--24677
"001101111100000000011111111111111001",--24678
"010011000011000000100000000000001000",--24679
"001101000000000000010000000100000000",--24680
"001101111100000000101111111111111010",--24681
"001101111100000000111111111111111011",--24682
"001001111100000111111111111111111000",--24683
"101001111100010111100000000000001001",--24684
"000111000000000000000100101110010000",--24685
"101001111100000111100000000000001001",--24686
"001101111100000111111111111111111000",--24687
"001101111100000000011111111111111001",--24688
"010011000011000000110000000000001000",--24689
"001101000000000000010000000100000001",--24690
"001101111100000000101111111111111010",--24691
"001101111100000000111111111111111011",--24692
"001001111100000111111111111111111000",--24693
"101001111100010111100000000000001001",--24694
"000111000000000000000100101110010000",--24695
"101001111100000111100000000000001001",--24696
"001101111100000111111111111111111000",--24697
"001101111100000000011111111111111001",--24698
"010011000011000001000000000000001000",--24699
"001101000000000000010000000100000010",--24700
"001101111100000000101111111111111010",--24701
"001101111100000000111111111111111011",--24702
"001001111100000111111111111111111000",--24703
"101001111100010111100000000000001001",--24704
"000111000000000000000100101110010000",--24705
"101001111100000111100000000000001001",--24706
"001101111100000111111111111111111000",--24707
"001101111100000000011111111111111101",--24708
"001101111100000000111111111111111100",--24709
"001100000110000000010001000000000000",--24710
"001111000000000000110000000100011101",--24711
"001111000100000001000000000000000000",--24712
"001111000000000001010000000100100000",--24713
"111110001000001001010010000000000000",--24714
"111110000110000001000001100000000000",--24715
"001011000000000000110000000100011101",--24716
"001111000000000000110000000100011110",--24717
"001111000100000001000000000000000001",--24718
"001111000000000001010000000100100001",--24719
"111110001000001001010010000000000000",--24720
"111110000110000001000001100000000000",--24721
"001011000000000000110000000100011110",--24722
"001111000000000000110000000100011111",--24723
"001111000100000001000000000000000010",--24724
"001111000000000001010000000100100010",--24725
"111110001000001001010010000000000000",--24726
"111110000110000001000001100000000000",--24727
"001011000000000000110000000100011111",--24728
"001101111100000000011111111111111101",--24729
"101001000010000000010000000000000001",--24730
"011011000010000001011111100000000000",--24731
"001101111100000000111111111111111110",--24732
"001100000110000000010001000000000000",--24733
"010111000100000000001111100000000000",--24734
"001101111100000001001111111111111111",--24735
"001100001000000000010001000000000000",--24736
"010000000101000000000000000000101101",--24737
"001101111100000000100000000000000000",--24738
"001101000100000001010000000000000101",--24739
"001101000100000001100000000000000111",--24740
"001101000100000001110000000000000001",--24741
"001101000100000010000000000000000100",--24742
"001100001010000000010010100000000000",--24743
"001111001010000000110000000000000000",--24744
"001011000000000000110000000100100000",--24745
"001111001010000000110000000000000001",--24746
"001011000000000000110000000100100001",--24747
"001111001010000000110000000000000010",--24748
"001011000000000000110000000100100010",--24749
"001101000100000001010000000000000110",--24750
"001101001010000001010000000000000000",--24751
"001100001100000000010001000000000000",--24752
"001100001110000000010001100000000000",--24753
"001001111100000010001111111111111100",--24754
"001001111100000000011111111111111011",--24755
"101000001011111000000000100000000000",--24756
"001001111100000111111111111111111010",--24757
"101001111100010111100000000000000111",--24758
"000111000000000000000101000111001101",--24759
"101001111100000111100000000000000111",--24760
"001101111100000111111111111111111010",--24761
"001101111100000000011111111111111011",--24762
"001101111100000000111111111111111100",--24763
"001100000110000000010001000000000000",--24764
"001111000000000000110000000100011101",--24765
"001111000100000001000000000000000000",--24766
"001111000000000001010000000100100000",--24767
"111110001000001001010010000000000000",--24768
"111110000110000001000001100000000000",--24769
"001011000000000000110000000100011101",--24770
"001111000000000000110000000100011110",--24771
"001111000100000001000000000000000001",--24772
"001111000000000001010000000100100001",--24773
"111110001000001001010010000000000000",--24774
"111110000110000001000001100000000000",--24775
"001011000000000000110000000100011110",--24776
"001111000000000000110000000100011111",--24777
"001111000100000001000000000000000010",--24778
"001111000000000001010000000100100010",--24779
"111110001000001001010010000000000000",--24780
"111110000110000001000001100000000000",--24781
"001011000000000000110000000100011111",--24782
"101001000010000000100000000000000001",--24783
"011011000100000001011111100000000000",--24784
"001101111100000000111111111111111110",--24785
"001100000110000000100000100000000000",--24786
"010111000010000000001111100000000000",--24787
"001101111100000000111111111111111111",--24788
"001100000110000000100000100000000000",--24789
"001001111100000000101111111111111100",--24790
"010000000011000000000000000000000110",--24791
"001101111100000000010000000000000000",--24792
"001001111100000111111111111111111011",--24793
"101001111100010111100000000000000110",--24794
"000111000000000000000101011001110000",--24795
"101001111100000111100000000000000110",--24796
"001101111100000111111111111111111011",--24797
"001101111100000000011111111111111100",--24798
"101001000010000000100000000000000001",--24799
"001101111100000000010000000000000000",--24800
"011011000100000001011111100000000000",--24801
"000101000000000000000101101010010001",--24802
"001101001110000001110000000000000011",--24803
"001100001110000001100011100000000000",--24804
"010000001111000000000000000001011100",--24805
"001100000110000000010011100000000000",--24806
"001101001110000001110000000000000101",--24807
"101001000010010010000000000000000001",--24808
"001100001000000010000100000000000000",--24809
"001101010000000010000000000000000101",--24810
"001100001000000000010100100000000000",--24811
"001101010010000010010000000000000101",--24812
"101001000010000010100000000000000001",--24813
"001100001000000010100101000000000000",--24814
"001101010100000010100000000000000101",--24815
"001100001010000000010101100000000000",--24816
"001101010110000010110000000000000101",--24817
"001100001110000001100011100000000000",--24818
"001111001110000000110000000000000000",--24819
"001011000000000000110000000100100000",--24820
"001111001110000000110000000000000001",--24821
"001011000000000000110000000100100001",--24822
"001111001110000000110000000000000010",--24823
"001011000000000000110000000100100010",--24824
"001100010000000001100011100000000000",--24825
"001111000000000000110000000100100000",--24826
"001111001110000001000000000000000000",--24827
"111110000110000001000001100000000000",--24828
"001011000000000000110000000100100000",--24829
"001111000000000000110000000100100001",--24830
"001111001110000001000000000000000001",--24831
"111110000110000001000001100000000000",--24832
"001011000000000000110000000100100001",--24833
"001111000000000000110000000100100010",--24834
"001111001110000001000000000000000010",--24835
"111110000110000001000001100000000000",--24836
"001011000000000000110000000100100010",--24837
"001100010010000001100011100000000000",--24838
"001111000000000000110000000100100000",--24839
"001111001110000001000000000000000000",--24840
"111110000110000001000001100000000000",--24841
"001011000000000000110000000100100000",--24842
"001111000000000000110000000100100001",--24843
"001111001110000001000000000000000001",--24844
"111110000110000001000001100000000000",--24845
"001011000000000000110000000100100001",--24846
"001111000000000000110000000100100010",--24847
"001111001110000001000000000000000010",--24848
"111110000110000001000001100000000000",--24849
"001011000000000000110000000100100010",--24850
"001100010100000001100011100000000000",--24851
"001111000000000000110000000100100000",--24852
"001111001110000001000000000000000000",--24853
"111110000110000001000001100000000000",--24854
"001011000000000000110000000100100000",--24855
"001111000000000000110000000100100001",--24856
"001111001110000001000000000000000001",--24857
"111110000110000001000001100000000000",--24858
"001011000000000000110000000100100001",--24859
"001111000000000000110000000100100010",--24860
"001111001110000001000000000000000010",--24861
"111110000110000001000001100000000000",--24862
"001011000000000000110000000100100010",--24863
"001100010110000001100011100000000000",--24864
"001111000000000000110000000100100000",--24865
"001111001110000001000000000000000000",--24866
"111110000110000001000001100000000000",--24867
"001011000000000000110000000100100000",--24868
"001111000000000000110000000100100001",--24869
"001111001110000001000000000000000001",--24870
"111110000110000001000001100000000000",--24871
"001011000000000000110000000100100001",--24872
"001111000000000000110000000100100010",--24873
"001111001110000001000000000000000010",--24874
"111110000110000001000001100000000000",--24875
"001011000000000000110000000100100010",--24876
"001100001000000000010011100000000000",--24877
"001101001110000001110000000000000100",--24878
"001100001110000001100011100000000000",--24879
"001111000000000000110000000100011101",--24880
"001111001110000001000000000000000000",--24881
"001111000000000001010000000100100000",--24882
"111110001000001001010010000000000000",--24883
"111110000110000001000001100000000000",--24884
"001011000000000000110000000100011101",--24885
"001111000000000000110000000100011110",--24886
"001111001110000001000000000000000001",--24887
"001111000000000001010000000100100001",--24888
"111110001000001001010010000000000000",--24889
"111110000110000001000001100000000000",--24890
"001011000000000000110000000100011110",--24891
"001111000000000000110000000100011111",--24892
"001111001110000001000000000000000010",--24893
"001111000000000001010000000100100010",--24894
"111110001000001001010010000000000000",--24895
"111110000110000001000001100000000000",--24896
"001011000000000000110000000100011111",--24897
"101001001100000001100000000000000001",--24898
"011011001100000001011111100000000000",--24899
"001100001000000000010011100000000000",--24900
"001101001110000010000000000000000010",--24901
"001100010000000001100100000000000000",--24902
"010111010000000000001111100000000000",--24903
"001100001000000000010100000000000000",--24904
"001101010000000010000000000000000010",--24905
"001100010000000001100100000000000000",--24906
"001100000110000000010100100000000000",--24907
"001101010010000010010000000000000010",--24908
"001100010010000001100100100000000000",--24909
"011100010011000010000000000000010100",--24910
"001100001010000000010100100000000000",--24911
"001101010010000010010000000000000010",--24912
"001100010010000001100100100000000000",--24913
"011100010011000010000000000000001110",--24914
"101001000010010010010000000000000001",--24915
"001100001000000010010100100000000000",--24916
"001101010010000010010000000000000010",--24917
"001100010010000001100100100000000000",--24918
"011100010011000010000000000000000111",--24919
"101001000010000010010000000000000001",--24920
"001100001000000010010100100000000000",--24921
"001101010010000010010000000000000010",--24922
"001100010010000001100100100000000000",--24923
"010000010011000010000000000001010001",--24924
"011011001100000001011111100000000000",--24925
"000101000000000000000110000101100100",--24926
"011011001100000001011111100000000000",--24927
"000101000000000000000110000101100100",--24928
"011011001100000001011111100000000000",--24929
"000101000000000000000110000101100100",--24930
"011011001100000001011111100000000000",--24931
"001100001000000000010000100000000000",--24932
"001101000010000000100000000000000010",--24933
"001100000100000001100001100000000000",--24934
"010111000110000000001111100000000000",--24935
"001101000010000000110000000000000011",--24936
"001100000110000001100010000000000000",--24937
"001001111100000000010000000000000000",--24938
"001001111100000000111111111111111111",--24939
"001001111100000000101111111111111110",--24940
"001001111100000001101111111111111101",--24941
"010000001001000000000000000000101010",--24942
"001101000010000001000000000000000101",--24943
"001101000010000001010000000000000111",--24944
"001101000010000001110000000000000001",--24945
"001101000010000010000000000000000100",--24946
"001100001000000001100010000000000000",--24947
"001111001000000000110000000000000000",--24948
"001011000000000000110000000100100000",--24949
"001111001000000000110000000000000001",--24950
"001011000000000000110000000100100001",--24951
"001111001000000000110000000000000010",--24952
"001011000000000000110000000100100010",--24953
"001101000010000001000000000000000110",--24954
"001101001000000000010000000000000000",--24955
"001100001010000001100001000000000000",--24956
"001100001110000001100001100000000000",--24957
"001001111100000010001111111111111100",--24958
"001001111100000111111111111111111011",--24959
"101001111100010111100000000000000110",--24960
"000111000000000000000101000111001101",--24961
"101001111100000111100000000000000110",--24962
"001101111100000111111111111111111011",--24963
"001101111100000000011111111111111101",--24964
"001101111100000000111111111111111100",--24965
"001100000110000000010001000000000000",--24966
"001111000000000000110000000100011101",--24967
"001111000100000001000000000000000000",--24968
"001111000000000001010000000100100000",--24969
"111110001000001001010010000000000000",--24970
"111110000110000001000001100000000000",--24971
"001011000000000000110000000100011101",--24972
"001111000000000000110000000100011110",--24973
"001111000100000001000000000000000001",--24974
"001111000000000001010000000100100001",--24975
"111110001000001001010010000000000000",--24976
"111110000110000001000001100000000000",--24977
"001011000000000000110000000100011110",--24978
"001111000000000000110000000100011111",--24979
"001111000100000001000000000000000010",--24980
"001111000000000001010000000100100010",--24981
"111110001000001001010010000000000000",--24982
"111110000110000001000001100000000000",--24983
"001011000000000000110000000100011111",--24984
"001101111100000000011111111111111101",--24985
"101001000010000000100000000000000001",--24986
"011011000100000001011111100000000000",--24987
"001101111100000000111111111111111110",--24988
"001100000110000000100000100000000000",--24989
"010111000010000000001111100000000000",--24990
"001101111100000000111111111111111111",--24991
"001100000110000000100000100000000000",--24992
"001001111100000000101111111111111100",--24993
"010000000011000000000000000000000110",--24994
"001101111100000000010000000000000000",--24995
"001001111100000111111111111111111011",--24996
"101001111100010111100000000000000110",--24997
"000111000000000000000101011001110000",--24998
"101001111100000111100000000000000110",--24999
"001101111100000111111111111111111011",--25000
"001101111100000000011111111111111100",--25001
"101001000010000000100000000000000001",--25002
"001101111100000000010000000000000000",--25003
"011011000100000001011111100000000000",--25004
"000101000000000000000101101010010001",--25005
"001101001110000001110000000000000011",--25006
"001100001110000001100011100000000000",--25007
"010000001111000000000000000001011100",--25008
"001100000110000000010011100000000000",--25009
"001101001110000001110000000000000101",--25010
"101001000010010010000000000000000001",--25011
"001100001000000010000100000000000000",--25012
"001101010000000010000000000000000101",--25013
"001100001000000000010100100000000000",--25014
"001101010010000010010000000000000101",--25015
"101001000010000010100000000000000001",--25016
"001100001000000010100101000000000000",--25017
"001101010100000010100000000000000101",--25018
"001100001010000000010101100000000000",--25019
"001101010110000010110000000000000101",--25020
"001100001110000001100011100000000000",--25021
"001111001110000000110000000000000000",--25022
"001011000000000000110000000100100000",--25023
"001111001110000000110000000000000001",--25024
"001011000000000000110000000100100001",--25025
"001111001110000000110000000000000010",--25026
"001011000000000000110000000100100010",--25027
"001100010000000001100011100000000000",--25028
"001111000000000000110000000100100000",--25029
"001111001110000001000000000000000000",--25030
"111110000110000001000001100000000000",--25031
"001011000000000000110000000100100000",--25032
"001111000000000000110000000100100001",--25033
"001111001110000001000000000000000001",--25034
"111110000110000001000001100000000000",--25035
"001011000000000000110000000100100001",--25036
"001111000000000000110000000100100010",--25037
"001111001110000001000000000000000010",--25038
"111110000110000001000001100000000000",--25039
"001011000000000000110000000100100010",--25040
"001100010010000001100011100000000000",--25041
"001111000000000000110000000100100000",--25042
"001111001110000001000000000000000000",--25043
"111110000110000001000001100000000000",--25044
"001011000000000000110000000100100000",--25045
"001111000000000000110000000100100001",--25046
"001111001110000001000000000000000001",--25047
"111110000110000001000001100000000000",--25048
"001011000000000000110000000100100001",--25049
"001111000000000000110000000100100010",--25050
"001111001110000001000000000000000010",--25051
"111110000110000001000001100000000000",--25052
"001011000000000000110000000100100010",--25053
"001100010100000001100011100000000000",--25054
"001111000000000000110000000100100000",--25055
"001111001110000001000000000000000000",--25056
"111110000110000001000001100000000000",--25057
"001011000000000000110000000100100000",--25058
"001111000000000000110000000100100001",--25059
"001111001110000001000000000000000001",--25060
"111110000110000001000001100000000000",--25061
"001011000000000000110000000100100001",--25062
"001111000000000000110000000100100010",--25063
"001111001110000001000000000000000010",--25064
"111110000110000001000001100000000000",--25065
"001011000000000000110000000100100010",--25066
"001100010110000001100011100000000000",--25067
"001111000000000000110000000100100000",--25068
"001111001110000001000000000000000000",--25069
"111110000110000001000001100000000000",--25070
"001011000000000000110000000100100000",--25071
"001111000000000000110000000100100001",--25072
"001111001110000001000000000000000001",--25073
"111110000110000001000001100000000000",--25074
"001011000000000000110000000100100001",--25075
"001111000000000000110000000100100010",--25076
"001111001110000001000000000000000010",--25077
"111110000110000001000001100000000000",--25078
"001011000000000000110000000100100010",--25079
"001100001000000000010011100000000000",--25080
"001101001110000001110000000000000100",--25081
"001100001110000001100011100000000000",--25082
"001111000000000000110000000100011101",--25083
"001111001110000001000000000000000000",--25084
"001111000000000001010000000100100000",--25085
"111110001000001001010010000000000000",--25086
"111110000110000001000001100000000000",--25087
"001011000000000000110000000100011101",--25088
"001111000000000000110000000100011110",--25089
"001111001110000001000000000000000001",--25090
"001111000000000001010000000100100001",--25091
"111110001000001001010010000000000000",--25092
"111110000110000001000001100000000000",--25093
"001011000000000000110000000100011110",--25094
"001111000000000000110000000100011111",--25095
"001111001110000001000000000000000010",--25096
"001111000000000001010000000100100010",--25097
"111110001000001001010010000000000000",--25098
"111110000110000001000001100000000000",--25099
"001011000000000000110000000100011111",--25100
"101001001100000001100000000000000001",--25101
"011011001100000001011111100000000000",--25102
"000101000000000000000110000000010101",--25103
"011011000100000001011111100000000000",--25104
"001101000010000000110000000000000010",--25105
"001100000110000000100010000000000000",--25106
"010111001000000000001111100000000000",--25107
"001101000010000001000000000000000011",--25108
"001100001000000000100010100000000000",--25109
"001001111100000001000000000000000000",--25110
"001001111100000000111111111111111111",--25111
"001001111100000000101111111111111110",--25112
"010000001011000000000000000100000001",--25113
"001101000010000001010000000000000110",--25114
"001101001010000001010000000000000000",--25115
"001011000000000000000000000100100000",--25116
"001011000000000000000000000100100001",--25117
"001011000000000000000000000100100010",--25118
"001101000010000001100000000000000111",--25119
"001101000010000001110000000000000001",--25120
"001101001010000001010000000011111110",--25121
"001100001100000000100011000000000000",--25122
"001100001110000000100011100000000000",--25123
"001111001110000000110000000000000000",--25124
"001011000000000000110000000100010010",--25125
"001111001110000000110000000000000001",--25126
"001011000000000000110000000100010011",--25127
"001111001110000000110000000000000010",--25128
"001011000000000000110000000100010100",--25129
"001101000000000010000000000110101010",--25130
"101001010000010010000000000000000001",--25131
"001001111100000000011111111111111101",--25132
"001001111100000001111111111111111100",--25133
"001001111100000001101111111111111011",--25134
"001001111100000001011111111111111010",--25135
"010111010001000000000000000011010111",--25136
"001101010000000010010000000101101101",--25137
"001101010010000010100000000000001010",--25138
"001101010010000010110000000000000001",--25139
"001111001110000000110000000000000000",--25140
"001101010010000011000000000000000101",--25141
"001111011000000001000000000000000000",--25142
"111110000110010001000001100000000000",--25143
"001011010100000000110000000000000000",--25144
"001111001110000000110000000000000001",--25145
"001111011000000001000000000000000001",--25146
"111110000110010001000001100000000000",--25147
"001011010100000000110000000000000001",--25148
"001111001110000000110000000000000010",--25149
"001111011000000001000000000000000010",--25150
"111110000110010001000001100000000000",--25151
"001011010100000000110000000000000010",--25152
"011111010111000000100000000000001110",--25153
"001101010010000010010000000000000100",--25154
"001111010100000000110000000000000000",--25155
"001111010100000001000000000000000001",--25156
"001111010100000001010000000000000010",--25157
"001111010010000001100000000000000000",--25158
"111110001100001000110001100000000000",--25159
"001111010010000001100000000000000001",--25160
"111110001100001001000010000000000000",--25161
"111110000110000001000001100000000000",--25162
"001111010010000001000000000000000010",--25163
"111110001000001001010010000000000000",--25164
"111110000110000001000001100000000000",--25165
"001011010100000000110000000000000011",--25166
"000101000000000000000110001001110101",--25167
"010111010111000000100000000000100100",--25168
"001111010100000000110000000000000000",--25169
"001111010100000001000000000000000001",--25170
"001111010100000001010000000000000010",--25171
"111110000110001000110011000000000000",--25172
"001101010010000011000000000000000100",--25173
"001111011000000001110000000000000000",--25174
"111110001100001001110011000000000000",--25175
"111110001000001001000011100000000000",--25176
"001111011000000010000000000000000001",--25177
"111110001110001010000011100000000000",--25178
"111110001100000001110011000000000000",--25179
"111110001010001001010011100000000000",--25180
"001111011000000010000000000000000010",--25181
"111110001110001010000011100000000000",--25182
"111110001100000001110011000000000000",--25183
"001101010010000011000000000000000011",--25184
"011100011001000000000000000000000011",--25185
"101110001101111000000001100000000000",--25186
"011111010111000000110000000000010000",--25187
"000101000000000000000110001001110011",--25188
"111110001000001001010011100000000000",--25189
"001101010010000010010000000000001001",--25190
"001111010010000010000000000000000000",--25191
"111110001110001010000011100000000000",--25192
"111110001100000001110011000000000000",--25193
"111110001010001000110010100000000000",--25194
"001111010010000001110000000000000001",--25195
"111110001010001001110010100000000000",--25196
"111110001100000001010010100000000000",--25197
"111110000110001001000001100000000000",--25198
"001111010010000001000000000000000010",--25199
"111110000110001001000001100000000000",--25200
"111110001010000000110001100000000000",--25201
"011111010111000000110000000000000001",--25202
"111110000110010000010001100000000000",--25203
"001011010100000000110000000000000011",--25204
"101001010000010010000000000000000001",--25205
"010111010001000000000000000010010001",--25206
"001101010000000010010000000101101101",--25207
"001101010010000010100000000000001010",--25208
"001101010010000010110000000000000001",--25209
"001111001110000000110000000000000000",--25210
"001101010010000011000000000000000101",--25211
"001111011000000001000000000000000000",--25212
"111110000110010001000001100000000000",--25213
"001011010100000000110000000000000000",--25214
"001111001110000000110000000000000001",--25215
"001111011000000001000000000000000001",--25216
"111110000110010001000001100000000000",--25217
"001011010100000000110000000000000001",--25218
"001111001110000000110000000000000010",--25219
"001111011000000001000000000000000010",--25220
"111110000110010001000001100000000000",--25221
"001011010100000000110000000000000010",--25222
"011111010111000000100000000000001110",--25223
"001101010010000010010000000000000100",--25224
"001111010100000000110000000000000000",--25225
"001111010100000001000000000000000001",--25226
"001111010100000001010000000000000010",--25227
"001111010010000001100000000000000000",--25228
"111110001100001000110001100000000000",--25229
"001111010010000001100000000000000001",--25230
"111110001100001001000010000000000000",--25231
"111110000110000001000001100000000000",--25232
"001111010010000001000000000000000010",--25233
"111110001000001001010010000000000000",--25234
"111110000110000001000001100000000000",--25235
"001011010100000000110000000000000011",--25236
"000101000000000000000110001010111011",--25237
"010111010111000000100000000000100100",--25238
"001111010100000000110000000000000000",--25239
"001111010100000001000000000000000001",--25240
"001111010100000001010000000000000010",--25241
"111110000110001000110011000000000000",--25242
"001101010010000011000000000000000100",--25243
"001111011000000001110000000000000000",--25244
"111110001100001001110011000000000000",--25245
"111110001000001001000011100000000000",--25246
"001111011000000010000000000000000001",--25247
"111110001110001010000011100000000000",--25248
"111110001100000001110011000000000000",--25249
"111110001010001001010011100000000000",--25250
"001111011000000010000000000000000010",--25251
"111110001110001010000011100000000000",--25252
"111110001100000001110011000000000000",--25253
"001101010010000011000000000000000011",--25254
"011100011001000000000000000000000011",--25255
"101110001101111000000001100000000000",--25256
"011111010111000000110000000000010000",--25257
"000101000000000000000110001010111001",--25258
"111110001000001001010011100000000000",--25259
"001101010010000010010000000000001001",--25260
"001111010010000010000000000000000000",--25261
"111110001110001010000011100000000000",--25262
"111110001100000001110011000000000000",--25263
"111110001010001000110010100000000000",--25264
"001111010010000001110000000000000001",--25265
"111110001010001001110010100000000000",--25266
"111110001100000001010010100000000000",--25267
"111110000110001001000001100000000000",--25268
"001111010010000001000000000000000010",--25269
"111110000110001001000001100000000000",--25270
"111110001010000000110001100000000000",--25271
"011111010111000000110000000000000001",--25272
"111110000110010000010001100000000000",--25273
"001011010100000000110000000000000011",--25274
"101001010000010010000000000000000001",--25275
"010111010001000000000000000001001011",--25276
"001101010000000010010000000101101101",--25277
"001101010010000010100000000000001010",--25278
"001101010010000010110000000000000001",--25279
"001111001110000000110000000000000000",--25280
"001101010010000011000000000000000101",--25281
"001111011000000001000000000000000000",--25282
"111110000110010001000001100000000000",--25283
"001011010100000000110000000000000000",--25284
"001111001110000000110000000000000001",--25285
"001111011000000001000000000000000001",--25286
"111110000110010001000001100000000000",--25287
"001011010100000000110000000000000001",--25288
"001111001110000000110000000000000010",--25289
"001111011000000001000000000000000010",--25290
"111110000110010001000001100000000000",--25291
"001011010100000000110000000000000010",--25292
"011111010111000000100000000000001110",--25293
"001101010010000010010000000000000100",--25294
"001111010100000000110000000000000000",--25295
"001111010100000001000000000000000001",--25296
"001111010100000001010000000000000010",--25297
"001111010010000001100000000000000000",--25298
"111110001100001000110001100000000000",--25299
"001111010010000001100000000000000001",--25300
"111110001100001001000010000000000000",--25301
"111110000110000001000001100000000000",--25302
"001111010010000001000000000000000010",--25303
"111110001000001001010010000000000000",--25304
"111110000110000001000001100000000000",--25305
"001011010100000000110000000000000011",--25306
"000101000000000000000110001100000001",--25307
"010111010111000000100000000000100100",--25308
"001111010100000000110000000000000000",--25309
"001111010100000001000000000000000001",--25310
"001111010100000001010000000000000010",--25311
"111110000110001000110011000000000000",--25312
"001101010010000011000000000000000100",--25313
"001111011000000001110000000000000000",--25314
"111110001100001001110011000000000000",--25315
"111110001000001001000011100000000000",--25316
"001111011000000010000000000000000001",--25317
"111110001110001010000011100000000000",--25318
"111110001100000001110011000000000000",--25319
"111110001010001001010011100000000000",--25320
"001111011000000010000000000000000010",--25321
"111110001110001010000011100000000000",--25322
"111110001100000001110011000000000000",--25323
"001101010010000011000000000000000011",--25324
"011100011001000000000000000000000011",--25325
"101110001101111000000001100000000000",--25326
"011111010111000000110000000000010000",--25327
"000101000000000000000110001011111111",--25328
"111110001000001001010011100000000000",--25329
"001101010010000010010000000000001001",--25330
"001111010010000010000000000000000000",--25331
"111110001110001010000011100000000000",--25332
"111110001100000001110011000000000000",--25333
"111110001010001000110010100000000000",--25334
"001111010010000001110000000000000001",--25335
"111110001010001001110010100000000000",--25336
"111110001100000001010010100000000000",--25337
"111110000110001001000001100000000000",--25338
"001111010010000001000000000000000010",--25339
"111110000110001001000001100000000000",--25340
"111110001010000000110001100000000000",--25341
"011111010111000000110000000000000001",--25342
"111110000110010000010001100000000000",--25343
"001011010100000000110000000000000011",--25344
"101001010000010000100000000000000001",--25345
"101000001111111000000000100000000000",--25346
"001001111100000111111111111111111001",--25347
"101001111100010111100000000000001000",--25348
"000111000000000000000000011001101110",--25349
"101001111100000111100000000000001000",--25350
"001101111100000111111111111111111001",--25351
"101001000000000001000000000001110110",--25352
"001101111100000000011111111111111010",--25353
"001101111100000000101111111111111011",--25354
"001101111100000000111111111111111100",--25355
"001001111100000111111111111111111001",--25356
"101001111100010111100000000000001000",--25357
"000111000000000000000100000011011010",--25358
"101001111100000111100000000000001000",--25359
"001101111100000111111111111111111001",--25360
"001101111100000000011111111111111101",--25361
"001101000010000000100000000000000101",--25362
"001101111100000000111111111111111110",--25363
"001100000100000000110001000000000000",--25364
"001111000000000000110000000100100000",--25365
"001011000100000000110000000000000000",--25366
"001111000000000000110000000100100001",--25367
"001011000100000000110000000000000001",--25368
"001111000000000000110000000100100010",--25369
"001011000100000000110000000000000010",--25370
"001101111100000000101111111111111110",--25371
"101001000100000000100000000000000001",--25372
"011011000100000001011111100000000000",--25373
"001101111100000001001111111111111111",--25374
"001100001000000000100001100000000000",--25375
"010111000110000000001111100000000000",--25376
"001101111100000001010000000000000000",--25377
"001100001010000000100001100000000000",--25378
"001001111100000000101111111111111101",--25379
"010000000111000000000000000011011110",--25380
"001101000010000000110000000000000110",--25381
"001101000110000000110000000000000000",--25382
"001011000000000000000000000100100000",--25383
"001011000000000000000000000100100001",--25384
"001011000000000000000000000100100010",--25385
"001101000010000001100000000000000111",--25386
"001101000010000001110000000000000001",--25387
"001101000110000000110000000011111110",--25388
"001100001100000000100011000000000000",--25389
"001100001110000000100011100000000000",--25390
"001111001110000000110000000000000000",--25391
"001011000000000000110000000100010010",--25392
"001111001110000000110000000000000001",--25393
"001011000000000000110000000100010011",--25394
"001111001110000000110000000000000010",--25395
"001011000000000000110000000100010100",--25396
"001101000000000010000000000110101010",--25397
"101001010000010010000000000000000001",--25398
"001001111100000000011111111111111100",--25399
"001001111100000001111111111111111011",--25400
"001001111100000001101111111111111010",--25401
"001001111100000000111111111111111001",--25402
"010111010001000000000000000010010001",--25403
"001101010000000010010000000101101101",--25404
"001101010010000010100000000000001010",--25405
"001101010010000010110000000000000001",--25406
"001111001110000000110000000000000000",--25407
"001101010010000011000000000000000101",--25408
"001111011000000001000000000000000000",--25409
"111110000110010001000001100000000000",--25410
"001011010100000000110000000000000000",--25411
"001111001110000000110000000000000001",--25412
"001111011000000001000000000000000001",--25413
"111110000110010001000001100000000000",--25414
"001011010100000000110000000000000001",--25415
"001111001110000000110000000000000010",--25416
"001111011000000001000000000000000010",--25417
"111110000110010001000001100000000000",--25418
"001011010100000000110000000000000010",--25419
"011111010111000000100000000000001110",--25420
"001101010010000010010000000000000100",--25421
"001111010100000000110000000000000000",--25422
"001111010100000001000000000000000001",--25423
"001111010100000001010000000000000010",--25424
"001111010010000001100000000000000000",--25425
"111110001100001000110001100000000000",--25426
"001111010010000001100000000000000001",--25427
"111110001100001001000010000000000000",--25428
"111110000110000001000001100000000000",--25429
"001111010010000001000000000000000010",--25430
"111110001000001001010010000000000000",--25431
"111110000110000001000001100000000000",--25432
"001011010100000000110000000000000011",--25433
"000101000000000000000110001110000000",--25434
"010111010111000000100000000000100100",--25435
"001111010100000000110000000000000000",--25436
"001111010100000001000000000000000001",--25437
"001111010100000001010000000000000010",--25438
"111110000110001000110011000000000000",--25439
"001101010010000011000000000000000100",--25440
"001111011000000001110000000000000000",--25441
"111110001100001001110011000000000000",--25442
"111110001000001001000011100000000000",--25443
"001111011000000010000000000000000001",--25444
"111110001110001010000011100000000000",--25445
"111110001100000001110011000000000000",--25446
"111110001010001001010011100000000000",--25447
"001111011000000010000000000000000010",--25448
"111110001110001010000011100000000000",--25449
"111110001100000001110011000000000000",--25450
"001101010010000011000000000000000011",--25451
"011100011001000000000000000000000011",--25452
"101110001101111000000001100000000000",--25453
"011111010111000000110000000000010000",--25454
"000101000000000000000110001101111110",--25455
"111110001000001001010011100000000000",--25456
"001101010010000010010000000000001001",--25457
"001111010010000010000000000000000000",--25458
"111110001110001010000011100000000000",--25459
"111110001100000001110011000000000000",--25460
"111110001010001000110010100000000000",--25461
"001111010010000001110000000000000001",--25462
"111110001010001001110010100000000000",--25463
"111110001100000001010010100000000000",--25464
"111110000110001001000001100000000000",--25465
"001111010010000001000000000000000010",--25466
"111110000110001001000001100000000000",--25467
"111110001010000000110001100000000000",--25468
"011111010111000000110000000000000001",--25469
"111110000110010000010001100000000000",--25470
"001011010100000000110000000000000011",--25471
"101001010000010010000000000000000001",--25472
"010111010001000000000000000001001011",--25473
"001101010000000010010000000101101101",--25474
"001101010010000010100000000000001010",--25475
"001101010010000010110000000000000001",--25476
"001111001110000000110000000000000000",--25477
"001101010010000011000000000000000101",--25478
"001111011000000001000000000000000000",--25479
"111110000110010001000001100000000000",--25480
"001011010100000000110000000000000000",--25481
"001111001110000000110000000000000001",--25482
"001111011000000001000000000000000001",--25483
"111110000110010001000001100000000000",--25484
"001011010100000000110000000000000001",--25485
"001111001110000000110000000000000010",--25486
"001111011000000001000000000000000010",--25487
"111110000110010001000001100000000000",--25488
"001011010100000000110000000000000010",--25489
"011111010111000000100000000000001110",--25490
"001101010010000010010000000000000100",--25491
"001111010100000000110000000000000000",--25492
"001111010100000001000000000000000001",--25493
"001111010100000001010000000000000010",--25494
"001111010010000001100000000000000000",--25495
"111110001100001000110001100000000000",--25496
"001111010010000001100000000000000001",--25497
"111110001100001001000010000000000000",--25498
"111110000110000001000001100000000000",--25499
"001111010010000001000000000000000010",--25500
"111110001000001001010010000000000000",--25501
"111110000110000001000001100000000000",--25502
"001011010100000000110000000000000011",--25503
"000101000000000000000110001111000110",--25504
"010111010111000000100000000000100100",--25505
"001111010100000000110000000000000000",--25506
"001111010100000001000000000000000001",--25507
"001111010100000001010000000000000010",--25508
"111110000110001000110011000000000000",--25509
"001101010010000011000000000000000100",--25510
"001111011000000001110000000000000000",--25511
"111110001100001001110011000000000000",--25512
"111110001000001001000011100000000000",--25513
"001111011000000010000000000000000001",--25514
"111110001110001010000011100000000000",--25515
"111110001100000001110011000000000000",--25516
"111110001010001001010011100000000000",--25517
"001111011000000010000000000000000010",--25518
"111110001110001010000011100000000000",--25519
"111110001100000001110011000000000000",--25520
"001101010010000011000000000000000011",--25521
"011100011001000000000000000000000011",--25522
"101110001101111000000001100000000000",--25523
"011111010111000000110000000000010000",--25524
"000101000000000000000110001111000100",--25525
"111110001000001001010011100000000000",--25526
"001101010010000010010000000000001001",--25527
"001111010010000010000000000000000000",--25528
"111110001110001010000011100000000000",--25529
"111110001100000001110011000000000000",--25530
"111110001010001000110010100000000000",--25531
"001111010010000001110000000000000001",--25532
"111110001010001001110010100000000000",--25533
"111110001100000001010010100000000000",--25534
"111110000110001001000001100000000000",--25535
"001111010010000001000000000000000010",--25536
"111110000110001001000001100000000000",--25537
"111110001010000000110001100000000000",--25538
"011111010111000000110000000000000001",--25539
"111110000110010000010001100000000000",--25540
"001011010100000000110000000000000011",--25541
"101001010000010000100000000000000001",--25542
"101000001111111000000000100000000000",--25543
"001001111100000111111111111111111000",--25544
"101001111100010111100000000000001001",--25545
"000111000000000000000000011001101110",--25546
"101001111100000111100000000000001001",--25547
"001101111100000111111111111111111000",--25548
"001101111100000000011111111111111001",--25549
"001101000010000000100000000001110110",--25550
"001101000100000000100000000000000000",--25551
"001111000100000000110000000000000000",--25552
"001101111100000000111111111111111010",--25553
"001111000110000001000000000000000000",--25554
"111110000110001001000001100000000000",--25555
"001111000100000001000000000000000001",--25556
"001111000110000001010000000000000001",--25557
"111110001000001001010010000000000000",--25558
"111110000110000001000001100000000000",--25559
"001111000100000001000000000000000010",--25560
"001111000110000001010000000000000010",--25561
"111110001000001001010010000000000000",--25562
"111110000110000001000001100000000000",--25563
"011010000111000000000000000000001010",--25564
"001101000010000000010000000001110111",--25565
"101111001001110001001011101111011010",--25566
"101111001001100001000111010000001101",--25567
"111110000110001001000001100000000000",--25568
"001001111100000111111111111111111000",--25569
"101001111100010111100000000000001001",--25570
"000111000000000000000011110001110100",--25571
"101001111100000111100000000000001001",--25572
"001101111100000111111111111111111000",--25573
"000101000000000000000110001111110000",--25574
"001101000010000000010000000001110110",--25575
"101111001001110001000011101111011010",--25576
"101111001001100001000111010000001101",--25577
"111110000110001001000001100000000000",--25578
"001001111100000111111111111111111000",--25579
"101001111100010111100000000000001001",--25580
"000111000000000000000011110001110100",--25581
"101001111100000111100000000000001001",--25582
"001101111100000111111111111111111000",--25583
"101001000000000001000000000001110100",--25584
"001101111100000000011111111111111001",--25585
"001101111100000000101111111111111010",--25586
"001101111100000000111111111111111011",--25587
"001001111100000111111111111111111000",--25588
"101001111100010111100000000000001001",--25589
"000111000000000000000100000011011010",--25590
"101001111100000111100000000000001001",--25591
"001101111100000111111111111111111000",--25592
"001101111100000000011111111111111100",--25593
"001101000010000000100000000000000101",--25594
"001101111100000000111111111111111101",--25595
"001100000100000000110001000000000000",--25596
"001111000000000000110000000100100000",--25597
"001011000100000000110000000000000000",--25598
"001111000000000000110000000100100001",--25599
"001011000100000000110000000000000001",--25600
"001111000000000000110000000100100010",--25601
"001011000100000000110000000000000010",--25602
"001101111100000000101111111111111101",--25603
"101001000100000000100000000000000001",--25604
"011011000100000001011111100000000000",--25605
"001101111100000001001111111111111111",--25606
"001100001000000000100001100000000000",--25607
"010111000110000000001111100000000000",--25608
"001101111100000001010000000000000000",--25609
"001100001010000000100001100000000000",--25610
"001001111100000000101111111111111100",--25611
"010000000111000000000000000100000001",--25612
"001101000010000000110000000000000110",--25613
"001101000110000000110000000000000000",--25614
"001011000000000000000000000100100000",--25615
"001011000000000000000000000100100001",--25616
"001011000000000000000000000100100010",--25617
"001101000010000001100000000000000111",--25618
"001101000010000001110000000000000001",--25619
"001101000110000000110000000011111110",--25620
"001100001100000000100011000000000000",--25621
"001100001110000000100011100000000000",--25622
"001111001110000000110000000000000000",--25623
"001011000000000000110000000100010010",--25624
"001111001110000000110000000000000001",--25625
"001011000000000000110000000100010011",--25626
"001111001110000000110000000000000010",--25627
"001011000000000000110000000100010100",--25628
"001101000000000010000000000110101010",--25629
"101001010000010010000000000000000001",--25630
"001001111100000000011111111111111011",--25631
"001001111100000001111111111111111010",--25632
"001001111100000001101111111111111001",--25633
"001001111100000000111111111111111000",--25634
"010111010001000000000000000011010111",--25635
"001101010000000010010000000101101101",--25636
"001101010010000010100000000000001010",--25637
"001101010010000010110000000000000001",--25638
"001111001110000000110000000000000000",--25639
"001101010010000011000000000000000101",--25640
"001111011000000001000000000000000000",--25641
"111110000110010001000001100000000000",--25642
"001011010100000000110000000000000000",--25643
"001111001110000000110000000000000001",--25644
"001111011000000001000000000000000001",--25645
"111110000110010001000001100000000000",--25646
"001011010100000000110000000000000001",--25647
"001111001110000000110000000000000010",--25648
"001111011000000001000000000000000010",--25649
"111110000110010001000001100000000000",--25650
"001011010100000000110000000000000010",--25651
"011111010111000000100000000000001110",--25652
"001101010010000010010000000000000100",--25653
"001111010100000000110000000000000000",--25654
"001111010100000001000000000000000001",--25655
"001111010100000001010000000000000010",--25656
"001111010010000001100000000000000000",--25657
"111110001100001000110001100000000000",--25658
"001111010010000001100000000000000001",--25659
"111110001100001001000010000000000000",--25660
"111110000110000001000001100000000000",--25661
"001111010010000001000000000000000010",--25662
"111110001000001001010010000000000000",--25663
"111110000110000001000001100000000000",--25664
"001011010100000000110000000000000011",--25665
"000101000000000000000110010001101000",--25666
"010111010111000000100000000000100100",--25667
"001111010100000000110000000000000000",--25668
"001111010100000001000000000000000001",--25669
"001111010100000001010000000000000010",--25670
"111110000110001000110011000000000000",--25671
"001101010010000011000000000000000100",--25672
"001111011000000001110000000000000000",--25673
"111110001100001001110011000000000000",--25674
"111110001000001001000011100000000000",--25675
"001111011000000010000000000000000001",--25676
"111110001110001010000011100000000000",--25677
"111110001100000001110011000000000000",--25678
"111110001010001001010011100000000000",--25679
"001111011000000010000000000000000010",--25680
"111110001110001010000011100000000000",--25681
"111110001100000001110011000000000000",--25682
"001101010010000011000000000000000011",--25683
"011100011001000000000000000000000011",--25684
"101110001101111000000001100000000000",--25685
"011111010111000000110000000000010000",--25686
"000101000000000000000110010001100110",--25687
"111110001000001001010011100000000000",--25688
"001101010010000010010000000000001001",--25689
"001111010010000010000000000000000000",--25690
"111110001110001010000011100000000000",--25691
"111110001100000001110011000000000000",--25692
"111110001010001000110010100000000000",--25693
"001111010010000001110000000000000001",--25694
"111110001010001001110010100000000000",--25695
"111110001100000001010010100000000000",--25696
"111110000110001001000001100000000000",--25697
"001111010010000001000000000000000010",--25698
"111110000110001001000001100000000000",--25699
"111110001010000000110001100000000000",--25700
"011111010111000000110000000000000001",--25701
"111110000110010000010001100000000000",--25702
"001011010100000000110000000000000011",--25703
"101001010000010010000000000000000001",--25704
"010111010001000000000000000010010001",--25705
"001101010000000010010000000101101101",--25706
"001101010010000010100000000000001010",--25707
"001101010010000010110000000000000001",--25708
"001111001110000000110000000000000000",--25709
"001101010010000011000000000000000101",--25710
"001111011000000001000000000000000000",--25711
"111110000110010001000001100000000000",--25712
"001011010100000000110000000000000000",--25713
"001111001110000000110000000000000001",--25714
"001111011000000001000000000000000001",--25715
"111110000110010001000001100000000000",--25716
"001011010100000000110000000000000001",--25717
"001111001110000000110000000000000010",--25718
"001111011000000001000000000000000010",--25719
"111110000110010001000001100000000000",--25720
"001011010100000000110000000000000010",--25721
"011111010111000000100000000000001110",--25722
"001101010010000010010000000000000100",--25723
"001111010100000000110000000000000000",--25724
"001111010100000001000000000000000001",--25725
"001111010100000001010000000000000010",--25726
"001111010010000001100000000000000000",--25727
"111110001100001000110001100000000000",--25728
"001111010010000001100000000000000001",--25729
"111110001100001001000010000000000000",--25730
"111110000110000001000001100000000000",--25731
"001111010010000001000000000000000010",--25732
"111110001000001001010010000000000000",--25733
"111110000110000001000001100000000000",--25734
"001011010100000000110000000000000011",--25735
"000101000000000000000110010010101110",--25736
"010111010111000000100000000000100100",--25737
"001111010100000000110000000000000000",--25738
"001111010100000001000000000000000001",--25739
"001111010100000001010000000000000010",--25740
"111110000110001000110011000000000000",--25741
"001101010010000011000000000000000100",--25742
"001111011000000001110000000000000000",--25743
"111110001100001001110011000000000000",--25744
"111110001000001001000011100000000000",--25745
"001111011000000010000000000000000001",--25746
"111110001110001010000011100000000000",--25747
"111110001100000001110011000000000000",--25748
"111110001010001001010011100000000000",--25749
"001111011000000010000000000000000010",--25750
"111110001110001010000011100000000000",--25751
"111110001100000001110011000000000000",--25752
"001101010010000011000000000000000011",--25753
"011100011001000000000000000000000011",--25754
"101110001101111000000001100000000000",--25755
"011111010111000000110000000000010000",--25756
"000101000000000000000110010010101100",--25757
"111110001000001001010011100000000000",--25758
"001101010010000010010000000000001001",--25759
"001111010010000010000000000000000000",--25760
"111110001110001010000011100000000000",--25761
"111110001100000001110011000000000000",--25762
"111110001010001000110010100000000000",--25763
"001111010010000001110000000000000001",--25764
"111110001010001001110010100000000000",--25765
"111110001100000001010010100000000000",--25766
"111110000110001001000001100000000000",--25767
"001111010010000001000000000000000010",--25768
"111110000110001001000001100000000000",--25769
"111110001010000000110001100000000000",--25770
"011111010111000000110000000000000001",--25771
"111110000110010000010001100000000000",--25772
"001011010100000000110000000000000011",--25773
"101001010000010010000000000000000001",--25774
"010111010001000000000000000001001011",--25775
"001101010000000010010000000101101101",--25776
"001101010010000010100000000000001010",--25777
"001101010010000010110000000000000001",--25778
"001111001110000000110000000000000000",--25779
"001101010010000011000000000000000101",--25780
"001111011000000001000000000000000000",--25781
"111110000110010001000001100000000000",--25782
"001011010100000000110000000000000000",--25783
"001111001110000000110000000000000001",--25784
"001111011000000001000000000000000001",--25785
"111110000110010001000001100000000000",--25786
"001011010100000000110000000000000001",--25787
"001111001110000000110000000000000010",--25788
"001111011000000001000000000000000010",--25789
"111110000110010001000001100000000000",--25790
"001011010100000000110000000000000010",--25791
"011111010111000000100000000000001110",--25792
"001101010010000010010000000000000100",--25793
"001111010100000000110000000000000000",--25794
"001111010100000001000000000000000001",--25795
"001111010100000001010000000000000010",--25796
"001111010010000001100000000000000000",--25797
"111110001100001000110001100000000000",--25798
"001111010010000001100000000000000001",--25799
"111110001100001001000010000000000000",--25800
"111110000110000001000001100000000000",--25801
"001111010010000001000000000000000010",--25802
"111110001000001001010010000000000000",--25803
"111110000110000001000001100000000000",--25804
"001011010100000000110000000000000011",--25805
"000101000000000000000110010011110100",--25806
"010111010111000000100000000000100100",--25807
"001111010100000000110000000000000000",--25808
"001111010100000001000000000000000001",--25809
"001111010100000001010000000000000010",--25810
"111110000110001000110011000000000000",--25811
"001101010010000011000000000000000100",--25812
"001111011000000001110000000000000000",--25813
"111110001100001001110011000000000000",--25814
"111110001000001001000011100000000000",--25815
"001111011000000010000000000000000001",--25816
"111110001110001010000011100000000000",--25817
"111110001100000001110011000000000000",--25818
"111110001010001001010011100000000000",--25819
"001111011000000010000000000000000010",--25820
"111110001110001010000011100000000000",--25821
"111110001100000001110011000000000000",--25822
"001101010010000011000000000000000011",--25823
"011100011001000000000000000000000011",--25824
"101110001101111000000001100000000000",--25825
"011111010111000000110000000000010000",--25826
"000101000000000000000110010011110010",--25827
"111110001000001001010011100000000000",--25828
"001101010010000010010000000000001001",--25829
"001111010010000010000000000000000000",--25830
"111110001110001010000011100000000000",--25831
"111110001100000001110011000000000000",--25832
"111110001010001000110010100000000000",--25833
"001111010010000001110000000000000001",--25834
"111110001010001001110010100000000000",--25835
"111110001100000001010010100000000000",--25836
"111110000110001001000001100000000000",--25837
"001111010010000001000000000000000010",--25838
"111110000110001001000001100000000000",--25839
"111110001010000000110001100000000000",--25840
"011111010111000000110000000000000001",--25841
"111110000110010000010001100000000000",--25842
"001011010100000000110000000000000011",--25843
"101001010000010000100000000000000001",--25844
"101000001111111000000000100000000000",--25845
"001001111100000111111111111111110111",--25846
"101001111100010111100000000000001010",--25847
"000111000000000000000000011001101110",--25848
"101001111100000111100000000000001010",--25849
"001101111100000111111111111111110111",--25850
"101001000000000001000000000001110110",--25851
"001101111100000000011111111111111000",--25852
"001101111100000000101111111111111001",--25853
"001101111100000000111111111111111010",--25854
"001001111100000111111111111111110111",--25855
"101001111100010111100000000000001010",--25856
"000111000000000000000100000011011010",--25857
"101001111100000111100000000000001010",--25858
"001101111100000111111111111111110111",--25859
"001101111100000000011111111111111011",--25860
"001101000010000000100000000000000101",--25861
"001101111100000000111111111111111100",--25862
"001100000100000000110001000000000000",--25863
"001111000000000000110000000100100000",--25864
"001011000100000000110000000000000000",--25865
"001111000000000000110000000100100001",--25866
"001011000100000000110000000000000001",--25867
"001111000000000000110000000100100010",--25868
"001011000100000000110000000000000010",--25869
"001101111100000000101111111111111100",--25870
"101001000100000000100000000000000001",--25871
"011011000100000001011111100000000000",--25872
"001101111100000001001111111111111111",--25873
"001100001000000000100001100000000000",--25874
"010111000110000000001111100000000000",--25875
"001101111100000001000000000000000000",--25876
"001100001000000000100001100000000000",--25877
"001001111100000000101111111111111011",--25878
"010000000111000000000000000000011101",--25879
"001101000010000000110000000000000110",--25880
"001101000110000000110000000000000000",--25881
"001011000000000000000000000100100000",--25882
"001011000000000000000000000100100001",--25883
"001011000000000000000000000100100010",--25884
"001101000010000001000000000000000111",--25885
"001101000010000001010000000000000001",--25886
"001101000110000000110000000011111110",--25887
"001100001000000000100010000000000000",--25888
"001100001010000000100010100000000000",--25889
"001001111100000000011111111111111010",--25890
"101000001001111000000001000000000000",--25891
"101000000111111000000000100000000000",--25892
"101000001011111000000001100000000000",--25893
"001001111100000111111111111111111001",--25894
"101001111100010111100000000000001000",--25895
"000111000000000000000100101110010000",--25896
"101001111100000111100000000000001000",--25897
"001101111100000111111111111111111001",--25898
"001101111100000000011111111111111010",--25899
"001101000010000000100000000000000101",--25900
"001101111100000000111111111111111011",--25901
"001100000100000000110001000000000000",--25902
"001111000000000000110000000100100000",--25903
"001011000100000000110000000000000000",--25904
"001111000000000000110000000100100001",--25905
"001011000100000000110000000000000001",--25906
"001111000000000000110000000100100010",--25907
"001011000100000000110000000000000010",--25908
"001101111100000000101111111111111011",--25909
"101001000100000000100000000000000001",--25910
"011011000100000001011111100000000000",--25911
"000101000000000000000110001000010001",--25912
"010111000100000000001111100000000000",--25913
"001111000000000001100000000100011000",--25914
"001101000000000001000000000100011001",--25915
"101000000100010001000010000000000000",--25916
"101010001001101000000011100000000000",--25917
"111110001100001001110011000000000000",--25918
"001111000000000001110000000100001111",--25919
"111110001100001001110011100000000000",--25920
"111110001110000000110011100000000000",--25921
"001011000000000001110000000100000110",--25922
"001111000000000001110000000100010000",--25923
"111110001100001001110011100000000000",--25924
"111110001110000001000011100000000000",--25925
"001011000000000001110000000100000111",--25926
"001111000000000001110000000100010001",--25927
"111110001100001001110011000000000000",--25928
"111110001100000001010011000000000000",--25929
"001011000000000001100000000100001000",--25930
"001111000000000001100000000100000110",--25931
"111110001100001001100011000000000000",--25932
"001111000000000001110000000100000111",--25933
"111110001110001001110011100000000000",--25934
"111110001100000001110011000000000000",--25935
"001111000000000001110000000100001000",--25936
"111110001110001001110011100000000000",--25937
"111110001100000001110011000000000000",--25938
"111110001100100000000011000000000000",--25939
"011110001101000000000000000000000010",--25940
"101110000011111000000011000000000000",--25941
"000101000000000000000110010101011000",--25942
"111110001100011000000011000000000000",--25943
"001111000000000001110000000100000110",--25944
"111110001110001001100011100000000000",--25945
"001011000000000001110000000100000110",--25946
"001111000000000001110000000100000111",--25947
"111110001110001001100011100000000000",--25948
"001011000000000001110000000100000111",--25949
"001111000000000001110000000100001000",--25950
"111110001110001001100011000000000000",--25951
"001011000000000001100000000100001000",--25952
"001011000000000000000000000100011101",--25953
"001011000000000000000000000100011110",--25954
"001011000000000000000000000100011111",--25955
"001111000000000001100000000101100111",--25956
"001011000000000001100000000100010101",--25957
"001111000000000001100000000101101000",--25958
"001011000000000001100000000100010110",--25959
"001111000000000001100000000101101001",--25960
"001011000000000001100000000100010111",--25961
"001100000010000000100010100000000000",--25962
"001011111100000001010000000000000000",--25963
"001011111100000001001111111111111111",--25964
"001011111100000000111111111111111110",--25965
"001001111100000000111111111111111101",--25966
"001001111100000000011111111111111100",--25967
"001001111100000000101111111111111011",--25968
"101000001011111000000001100000000000",--25969
"101001000000000000100000000100000110",--25970
"101000000001111000000000100000000000",--25971
"101110000001111000000010000000000000",--25972
"101110000011111000000001100000000000",--25973
"001001111100000111111111111111111010",--25974
"101001111100010111100000000000000111",--25975
"000111000000000000000011010111001111",--25976
"101001111100000111100000000000000111",--25977
"001101111100000111111111111111111010",--25978
"001101111100000000011111111111111011",--25979
"001101111100000000111111111111111100",--25980
"001100000110000000010001000000000000",--25981
"001101000100000000100000000000000000",--25982
"001111000000000000110000000100011101",--25983
"001011000100000000110000000000000000",--25984
"001111000000000000110000000100011110",--25985
"001011000100000000110000000000000001",--25986
"001111000000000000110000000100011111",--25987
"001011000100000000110000000000000010",--25988
"001100000110000000010001000000000000",--25989
"001101000100000000100000000000000110",--25990
"001101111100000001001111111111111101",--25991
"001001000100000001000000000000000000",--25992
"001100000110000000010001000000000000",--25993
"001101000100000001010000000000000010",--25994
"001101001010000001100000000000000000",--25995
"010111001101000000000000001000001110",--25996
"001101000100000001100000000000000011",--25997
"001101001100000001110000000000000000",--25998
"001001111100000000101111111111111010",--25999
"001001111100000001101111111111111001",--26000
"001001111100000001011111111111111000",--26001
"010000001111000000000000000011011100",--26002
"001101000100000001110000000000000110",--26003
"001101001110000001110000000000000000",--26004
"001011000000000000000000000100100000",--26005
"001011000000000000000000000100100001",--26006
"001011000000000000000000000100100010",--26007
"001101000100000010000000000000000111",--26008
"001101000100000010010000000000000001",--26009
"001101001110000001110000000011111110",--26010
"001101010000000010000000000000000000",--26011
"001101010010000010010000000000000000",--26012
"001111010010000000110000000000000000",--26013
"001011000000000000110000000100010010",--26014
"001111010010000000110000000000000001",--26015
"001011000000000000110000000100010011",--26016
"001111010010000000110000000000000010",--26017
"001011000000000000110000000100010100",--26018
"001101000000000010100000000110101010",--26019
"101001010100010010100000000000000001",--26020
"001001111100000010011111111111110111",--26021
"001001111100000010001111111111110110",--26022
"001001111100000001111111111111110101",--26023
"010111010101000000000000000010010001",--26024
"001101010100000010110000000101101101",--26025
"001101010110000011000000000000001010",--26026
"001101010110000011010000000000000001",--26027
"001111010010000000110000000000000000",--26028
"001101010110000011100000000000000101",--26029
"001111011100000001000000000000000000",--26030
"111110000110010001000001100000000000",--26031
"001011011000000000110000000000000000",--26032
"001111010010000000110000000000000001",--26033
"001111011100000001000000000000000001",--26034
"111110000110010001000001100000000000",--26035
"001011011000000000110000000000000001",--26036
"001111010010000000110000000000000010",--26037
"001111011100000001000000000000000010",--26038
"111110000110010001000001100000000000",--26039
"001011011000000000110000000000000010",--26040
"011111011011000000100000000000001110",--26041
"001101010110000010110000000000000100",--26042
"001111011000000000110000000000000000",--26043
"001111011000000001000000000000000001",--26044
"001111011000000001010000000000000010",--26045
"001111010110000001100000000000000000",--26046
"111110001100001000110001100000000000",--26047
"001111010110000001100000000000000001",--26048
"111110001100001001000010000000000000",--26049
"111110000110000001000001100000000000",--26050
"001111010110000001000000000000000010",--26051
"111110001000001001010010000000000000",--26052
"111110000110000001000001100000000000",--26053
"001011011000000000110000000000000011",--26054
"000101000000000000000110010111101101",--26055
"010111011011000000100000000000100100",--26056
"001111011000000000110000000000000000",--26057
"001111011000000001000000000000000001",--26058
"001111011000000001010000000000000010",--26059
"111110000110001000110011000000000000",--26060
"001101010110000011100000000000000100",--26061
"001111011100000001110000000000000000",--26062
"111110001100001001110011000000000000",--26063
"111110001000001001000011100000000000",--26064
"001111011100000010000000000000000001",--26065
"111110001110001010000011100000000000",--26066
"111110001100000001110011000000000000",--26067
"111110001010001001010011100000000000",--26068
"001111011100000010000000000000000010",--26069
"111110001110001010000011100000000000",--26070
"111110001100000001110011000000000000",--26071
"001101010110000011100000000000000011",--26072
"011100011101000000000000000000000011",--26073
"101110001101111000000001100000000000",--26074
"011111011011000000110000000000010000",--26075
"000101000000000000000110010111101011",--26076
"111110001000001001010011100000000000",--26077
"001101010110000010110000000000001001",--26078
"001111010110000010000000000000000000",--26079
"111110001110001010000011100000000000",--26080
"111110001100000001110011000000000000",--26081
"111110001010001000110010100000000000",--26082
"001111010110000001110000000000000001",--26083
"111110001010001001110010100000000000",--26084
"111110001100000001010010100000000000",--26085
"111110000110001001000001100000000000",--26086
"001111010110000001000000000000000010",--26087
"111110000110001001000001100000000000",--26088
"111110001010000000110001100000000000",--26089
"011111011011000000110000000000000001",--26090
"111110000110010000010001100000000000",--26091
"001011011000000000110000000000000011",--26092
"101001010100010010100000000000000001",--26093
"010111010101000000000000000001001011",--26094
"001101010100000010110000000101101101",--26095
"001101010110000011000000000000001010",--26096
"001101010110000011010000000000000001",--26097
"001111010010000000110000000000000000",--26098
"001101010110000011100000000000000101",--26099
"001111011100000001000000000000000000",--26100
"111110000110010001000001100000000000",--26101
"001011011000000000110000000000000000",--26102
"001111010010000000110000000000000001",--26103
"001111011100000001000000000000000001",--26104
"111110000110010001000001100000000000",--26105
"001011011000000000110000000000000001",--26106
"001111010010000000110000000000000010",--26107
"001111011100000001000000000000000010",--26108
"111110000110010001000001100000000000",--26109
"001011011000000000110000000000000010",--26110
"011111011011000000100000000000001110",--26111
"001101010110000010110000000000000100",--26112
"001111011000000000110000000000000000",--26113
"001111011000000001000000000000000001",--26114
"001111011000000001010000000000000010",--26115
"001111010110000001100000000000000000",--26116
"111110001100001000110001100000000000",--26117
"001111010110000001100000000000000001",--26118
"111110001100001001000010000000000000",--26119
"111110000110000001000001100000000000",--26120
"001111010110000001000000000000000010",--26121
"111110001000001001010010000000000000",--26122
"111110000110000001000001100000000000",--26123
"001011011000000000110000000000000011",--26124
"000101000000000000000110011000110011",--26125
"010111011011000000100000000000100100",--26126
"001111011000000000110000000000000000",--26127
"001111011000000001000000000000000001",--26128
"001111011000000001010000000000000010",--26129
"111110000110001000110011000000000000",--26130
"001101010110000011100000000000000100",--26131
"001111011100000001110000000000000000",--26132
"111110001100001001110011000000000000",--26133
"111110001000001001000011100000000000",--26134
"001111011100000010000000000000000001",--26135
"111110001110001010000011100000000000",--26136
"111110001100000001110011000000000000",--26137
"111110001010001001010011100000000000",--26138
"001111011100000010000000000000000010",--26139
"111110001110001010000011100000000000",--26140
"111110001100000001110011000000000000",--26141
"001101010110000011100000000000000011",--26142
"011100011101000000000000000000000011",--26143
"101110001101111000000001100000000000",--26144
"011111011011000000110000000000010000",--26145
"000101000000000000000110011000110001",--26146
"111110001000001001010011100000000000",--26147
"001101010110000010110000000000001001",--26148
"001111010110000010000000000000000000",--26149
"111110001110001010000011100000000000",--26150
"111110001100000001110011000000000000",--26151
"111110001010001000110010100000000000",--26152
"001111010110000001110000000000000001",--26153
"111110001010001001110010100000000000",--26154
"111110001100000001010010100000000000",--26155
"111110000110001001000001100000000000",--26156
"001111010110000001000000000000000010",--26157
"111110000110001001000001100000000000",--26158
"111110001010000000110001100000000000",--26159
"011111011011000000110000000000000001",--26160
"111110000110010000010001100000000000",--26161
"001011011000000000110000000000000011",--26162
"101001010100010000100000000000000001",--26163
"101000010011111000000000100000000000",--26164
"001001111100000111111111111111110100",--26165
"101001111100010111100000000000001101",--26166
"000111000000000000000000011001101110",--26167
"101001111100000111100000000000001101",--26168
"001101111100000111111111111111110100",--26169
"001101111100000000011111111111110101",--26170
"001101000010000000100000000001110110",--26171
"001101000100000000100000000000000000",--26172
"001111000100000000110000000000000000",--26173
"001101111100000000111111111111110110",--26174
"001111000110000001000000000000000000",--26175
"111110000110001001000001100000000000",--26176
"001111000100000001000000000000000001",--26177
"001111000110000001010000000000000001",--26178
"111110001000001001010010000000000000",--26179
"111110000110000001000001100000000000",--26180
"001111000100000001000000000000000010",--26181
"001111000110000001010000000000000010",--26182
"111110001000001001010010000000000000",--26183
"111110000110000001000001100000000000",--26184
"011010000111000000000000000000001010",--26185
"001101000010000000010000000001110111",--26186
"101111001001110001001011101111011010",--26187
"101111001001100001000111010000001101",--26188
"111110000110001001000001100000000000",--26189
"001001111100000111111111111111110100",--26190
"101001111100010111100000000000001101",--26191
"000111000000000000000011110001110100",--26192
"101001111100000111100000000000001101",--26193
"001101111100000111111111111111110100",--26194
"000101000000000000000110011001011101",--26195
"001101000010000000010000000001110110",--26196
"101111001001110001000011101111011010",--26197
"101111001001100001000111010000001101",--26198
"111110000110001001000001100000000000",--26199
"001001111100000111111111111111110100",--26200
"101001111100010111100000000000001101",--26201
"000111000000000000000011110001110100",--26202
"101001111100000111100000000000001101",--26203
"001101111100000111111111111111110100",--26204
"101001000000000001000000000001110100",--26205
"001101111100000000011111111111110101",--26206
"001101111100000000101111111111110110",--26207
"001101111100000000111111111111110111",--26208
"001001111100000111111111111111110100",--26209
"101001111100010111100000000000001101",--26210
"000111000000000000000100000011011010",--26211
"101001111100000111100000000000001101",--26212
"001101111100000111111111111111110100",--26213
"001101111100000000011111111111111010",--26214
"001101000010000000100000000000000101",--26215
"001101000100000000100000000000000000",--26216
"001111000000000000110000000100100000",--26217
"001011000100000000110000000000000000",--26218
"001111000000000000110000000100100001",--26219
"001011000100000000110000000000000001",--26220
"001111000000000000110000000100100010",--26221
"001011000100000000110000000000000010",--26222
"001101111100000000011111111111111000",--26223
"001101000010000000100000000000000001",--26224
"010111000101000000000000000100101001",--26225
"001101111100000000101111111111111001",--26226
"001101000100000000110000000000000001",--26227
"010000000111000000000000000100000000",--26228
"001101111100000000111111111111111010",--26229
"001101000110000001000000000000000110",--26230
"001101001000000001000000000000000000",--26231
"001011000000000000000000000100100000",--26232
"001011000000000000000000000100100001",--26233
"001011000000000000000000000100100010",--26234
"001101000110000001010000000000000111",--26235
"001101000110000001100000000000000001",--26236
"001101001000000001000000000011111110",--26237
"001101001010000001010000000000000001",--26238
"001101001100000001100000000000000001",--26239
"001111001100000000110000000000000000",--26240
"001011000000000000110000000100010010",--26241
"001111001100000000110000000000000001",--26242
"001011000000000000110000000100010011",--26243
"001111001100000000110000000000000010",--26244
"001011000000000000110000000100010100",--26245
"001101000000000001110000000110101010",--26246
"101001001110010001110000000000000001",--26247
"001001111100000001101111111111110111",--26248
"001001111100000001011111111111110110",--26249
"001001111100000001001111111111110101",--26250
"010111001111000000000000000011010111",--26251
"001101001110000010000000000101101101",--26252
"001101010000000010010000000000001010",--26253
"001101010000000010100000000000000001",--26254
"001111001100000000110000000000000000",--26255
"001101010000000010110000000000000101",--26256
"001111010110000001000000000000000000",--26257
"111110000110010001000001100000000000",--26258
"001011010010000000110000000000000000",--26259
"001111001100000000110000000000000001",--26260
"001111010110000001000000000000000001",--26261
"111110000110010001000001100000000000",--26262
"001011010010000000110000000000000001",--26263
"001111001100000000110000000000000010",--26264
"001111010110000001000000000000000010",--26265
"111110000110010001000001100000000000",--26266
"001011010010000000110000000000000010",--26267
"011111010101000000100000000000001110",--26268
"001101010000000010000000000000000100",--26269
"001111010010000000110000000000000000",--26270
"001111010010000001000000000000000001",--26271
"001111010010000001010000000000000010",--26272
"001111010000000001100000000000000000",--26273
"111110001100001000110001100000000000",--26274
"001111010000000001100000000000000001",--26275
"111110001100001001000010000000000000",--26276
"111110000110000001000001100000000000",--26277
"001111010000000001000000000000000010",--26278
"111110001000001001010010000000000000",--26279
"111110000110000001000001100000000000",--26280
"001011010010000000110000000000000011",--26281
"000101000000000000000110011011010000",--26282
"010111010101000000100000000000100100",--26283
"001111010010000000110000000000000000",--26284
"001111010010000001000000000000000001",--26285
"001111010010000001010000000000000010",--26286
"111110000110001000110011000000000000",--26287
"001101010000000010110000000000000100",--26288
"001111010110000001110000000000000000",--26289
"111110001100001001110011000000000000",--26290
"111110001000001001000011100000000000",--26291
"001111010110000010000000000000000001",--26292
"111110001110001010000011100000000000",--26293
"111110001100000001110011000000000000",--26294
"111110001010001001010011100000000000",--26295
"001111010110000010000000000000000010",--26296
"111110001110001010000011100000000000",--26297
"111110001100000001110011000000000000",--26298
"001101010000000010110000000000000011",--26299
"011100010111000000000000000000000011",--26300
"101110001101111000000001100000000000",--26301
"011111010101000000110000000000010000",--26302
"000101000000000000000110011011001110",--26303
"111110001000001001010011100000000000",--26304
"001101010000000010000000000000001001",--26305
"001111010000000010000000000000000000",--26306
"111110001110001010000011100000000000",--26307
"111110001100000001110011000000000000",--26308
"111110001010001000110010100000000000",--26309
"001111010000000001110000000000000001",--26310
"111110001010001001110010100000000000",--26311
"111110001100000001010010100000000000",--26312
"111110000110001001000001100000000000",--26313
"001111010000000001000000000000000010",--26314
"111110000110001001000001100000000000",--26315
"111110001010000000110001100000000000",--26316
"011111010101000000110000000000000001",--26317
"111110000110010000010001100000000000",--26318
"001011010010000000110000000000000011",--26319
"101001001110010001110000000000000001",--26320
"010111001111000000000000000010010001",--26321
"001101001110000010000000000101101101",--26322
"001101010000000010010000000000001010",--26323
"001101010000000010100000000000000001",--26324
"001111001100000000110000000000000000",--26325
"001101010000000010110000000000000101",--26326
"001111010110000001000000000000000000",--26327
"111110000110010001000001100000000000",--26328
"001011010010000000110000000000000000",--26329
"001111001100000000110000000000000001",--26330
"001111010110000001000000000000000001",--26331
"111110000110010001000001100000000000",--26332
"001011010010000000110000000000000001",--26333
"001111001100000000110000000000000010",--26334
"001111010110000001000000000000000010",--26335
"111110000110010001000001100000000000",--26336
"001011010010000000110000000000000010",--26337
"011111010101000000100000000000001110",--26338
"001101010000000010000000000000000100",--26339
"001111010010000000110000000000000000",--26340
"001111010010000001000000000000000001",--26341
"001111010010000001010000000000000010",--26342
"001111010000000001100000000000000000",--26343
"111110001100001000110001100000000000",--26344
"001111010000000001100000000000000001",--26345
"111110001100001001000010000000000000",--26346
"111110000110000001000001100000000000",--26347
"001111010000000001000000000000000010",--26348
"111110001000001001010010000000000000",--26349
"111110000110000001000001100000000000",--26350
"001011010010000000110000000000000011",--26351
"000101000000000000000110011100010110",--26352
"010111010101000000100000000000100100",--26353
"001111010010000000110000000000000000",--26354
"001111010010000001000000000000000001",--26355
"001111010010000001010000000000000010",--26356
"111110000110001000110011000000000000",--26357
"001101010000000010110000000000000100",--26358
"001111010110000001110000000000000000",--26359
"111110001100001001110011000000000000",--26360
"111110001000001001000011100000000000",--26361
"001111010110000010000000000000000001",--26362
"111110001110001010000011100000000000",--26363
"111110001100000001110011000000000000",--26364
"111110001010001001010011100000000000",--26365
"001111010110000010000000000000000010",--26366
"111110001110001010000011100000000000",--26367
"111110001100000001110011000000000000",--26368
"001101010000000010110000000000000011",--26369
"011100010111000000000000000000000011",--26370
"101110001101111000000001100000000000",--26371
"011111010101000000110000000000010000",--26372
"000101000000000000000110011100010100",--26373
"111110001000001001010011100000000000",--26374
"001101010000000010000000000000001001",--26375
"001111010000000010000000000000000000",--26376
"111110001110001010000011100000000000",--26377
"111110001100000001110011000000000000",--26378
"111110001010001000110010100000000000",--26379
"001111010000000001110000000000000001",--26380
"111110001010001001110010100000000000",--26381
"111110001100000001010010100000000000",--26382
"111110000110001001000001100000000000",--26383
"001111010000000001000000000000000010",--26384
"111110000110001001000001100000000000",--26385
"111110001010000000110001100000000000",--26386
"011111010101000000110000000000000001",--26387
"111110000110010000010001100000000000",--26388
"001011010010000000110000000000000011",--26389
"101001001110010001110000000000000001",--26390
"010111001111000000000000000001001011",--26391
"001101001110000010000000000101101101",--26392
"001101010000000010010000000000001010",--26393
"001101010000000010100000000000000001",--26394
"001111001100000000110000000000000000",--26395
"001101010000000010110000000000000101",--26396
"001111010110000001000000000000000000",--26397
"111110000110010001000001100000000000",--26398
"001011010010000000110000000000000000",--26399
"001111001100000000110000000000000001",--26400
"001111010110000001000000000000000001",--26401
"111110000110010001000001100000000000",--26402
"001011010010000000110000000000000001",--26403
"001111001100000000110000000000000010",--26404
"001111010110000001000000000000000010",--26405
"111110000110010001000001100000000000",--26406
"001011010010000000110000000000000010",--26407
"011111010101000000100000000000001110",--26408
"001101010000000010000000000000000100",--26409
"001111010010000000110000000000000000",--26410
"001111010010000001000000000000000001",--26411
"001111010010000001010000000000000010",--26412
"001111010000000001100000000000000000",--26413
"111110001100001000110001100000000000",--26414
"001111010000000001100000000000000001",--26415
"111110001100001001000010000000000000",--26416
"111110000110000001000001100000000000",--26417
"001111010000000001000000000000000010",--26418
"111110001000001001010010000000000000",--26419
"111110000110000001000001100000000000",--26420
"001011010010000000110000000000000011",--26421
"000101000000000000000110011101011100",--26422
"010111010101000000100000000000100100",--26423
"001111010010000000110000000000000000",--26424
"001111010010000001000000000000000001",--26425
"001111010010000001010000000000000010",--26426
"111110000110001000110011000000000000",--26427
"001101010000000010110000000000000100",--26428
"001111010110000001110000000000000000",--26429
"111110001100001001110011000000000000",--26430
"111110001000001001000011100000000000",--26431
"001111010110000010000000000000000001",--26432
"111110001110001010000011100000000000",--26433
"111110001100000001110011000000000000",--26434
"111110001010001001010011100000000000",--26435
"001111010110000010000000000000000010",--26436
"111110001110001010000011100000000000",--26437
"111110001100000001110011000000000000",--26438
"001101010000000010110000000000000011",--26439
"011100010111000000000000000000000011",--26440
"101110001101111000000001100000000000",--26441
"011111010101000000110000000000010000",--26442
"000101000000000000000110011101011010",--26443
"111110001000001001010011100000000000",--26444
"001101010000000010000000000000001001",--26445
"001111010000000010000000000000000000",--26446
"111110001110001010000011100000000000",--26447
"111110001100000001110011000000000000",--26448
"111110001010001000110010100000000000",--26449
"001111010000000001110000000000000001",--26450
"111110001010001001110010100000000000",--26451
"111110001100000001010010100000000000",--26452
"111110000110001001000001100000000000",--26453
"001111010000000001000000000000000010",--26454
"111110000110001001000001100000000000",--26455
"111110001010000000110001100000000000",--26456
"011111010101000000110000000000000001",--26457
"111110000110010000010001100000000000",--26458
"001011010010000000110000000000000011",--26459
"101001001110010000100000000000000001",--26460
"101000001101111000000000100000000000",--26461
"001001111100000111111111111111110100",--26462
"101001111100010111100000000000001101",--26463
"000111000000000000000000011001101110",--26464
"101001111100000111100000000000001101",--26465
"001101111100000111111111111111110100",--26466
"101001000000000001000000000001110110",--26467
"001101111100000000011111111111110101",--26468
"001101111100000000101111111111110110",--26469
"001101111100000000111111111111110111",--26470
"001001111100000111111111111111110100",--26471
"101001111100010111100000000000001101",--26472
"000111000000000000000100000011011010",--26473
"101001111100000111100000000000001101",--26474
"001101111100000111111111111111110100",--26475
"001101111100000000011111111111111010",--26476
"001101000010000000100000000000000101",--26477
"001101000100000000100000000000000001",--26478
"001111000000000000110000000100100000",--26479
"001011000100000000110000000000000000",--26480
"001111000000000000110000000100100001",--26481
"001011000100000000110000000000000001",--26482
"001111000000000000110000000100100010",--26483
"001011000100000000110000000000000010",--26484
"001101111100000000011111111111111000",--26485
"001101000010000000010000000000000010",--26486
"010111000011000000000000000000100011",--26487
"001101111100000000011111111111111001",--26488
"001101000010000000010000000000000010",--26489
"010000000011000000000000000000011001",--26490
"001101111100000000011111111111111010",--26491
"001101000010000000100000000000000110",--26492
"001101000100000000100000000000000000",--26493
"001011000000000000000000000100100000",--26494
"001011000000000000000000000100100001",--26495
"001011000000000000000000000100100010",--26496
"001101000010000000110000000000000111",--26497
"001101000010000001000000000000000001",--26498
"001101000100000000010000000011111110",--26499
"001101000110000000100000000000000010",--26500
"001101001000000000110000000000000010",--26501
"001001111100000111111111111111110111",--26502
"101001111100010111100000000000001010",--26503
"000111000000000000000100101110010000",--26504
"101001111100000111100000000000001010",--26505
"001101111100000111111111111111110111",--26506
"001101111100000000011111111111111010",--26507
"001101000010000000100000000000000101",--26508
"001101000100000000100000000000000010",--26509
"001111000000000000110000000100100000",--26510
"001011000100000000110000000000000000",--26511
"001111000000000000110000000100100001",--26512
"001011000100000000110000000000000001",--26513
"001111000000000000110000000100100010",--26514
"001011000100000000110000000000000010",--26515
"101001000000000000100000000000000011",--26516
"001101111100000000011111111111111010",--26517
"001001111100000111111111111111110111",--26518
"101001111100010111100000000000001010",--26519
"000111000000000000000110001000010000",--26520
"101001111100000111100000000000001010",--26521
"001101111100000111111111111111110111",--26522
"001101111100000000011111111111111011",--26523
"101001000010010000010000000000000001",--26524
"010111000010000000001111100000000000",--26525
"001101111100000000101111111111111101",--26526
"101001000100000000100000000000000001",--26527
"010111000101000001000000000000000001",--26528
"101001000100010000100000000000000101",--26529
"001111000000000000110000000100011000",--26530
"001101000000000000110000000100011001",--26531
"101000000010010000110001100000000000",--26532
"101010000111101000000010000000000000",--26533
"111110000110001001000001100000000000",--26534
"001111000000000001000000000100001111",--26535
"111110000110001001000010000000000000",--26536
"001111111100000001011111111111111110",--26537
"111110001000000001010010000000000000",--26538
"001011000000000001000000000100000110",--26539
"001111000000000001000000000100010000",--26540
"111110000110001001000010000000000000",--26541
"001111111100000001101111111111111111",--26542
"111110001000000001100010000000000000",--26543
"001011000000000001000000000100000111",--26544
"001111000000000001000000000100010001",--26545
"111110000110001001000001100000000000",--26546
"001111111100000001000000000000000000",--26547
"111110000110000001000001100000000000",--26548
"001011000000000000110000000100001000",--26549
"001111000000000000110000000100000110",--26550
"111110000110001000110001100000000000",--26551
"001111000000000001110000000100000111",--26552
"111110001110001001110011100000000000",--26553
"111110000110000001110001100000000000",--26554
"001111000000000001110000000100001000",--26555
"111110001110001001110011100000000000",--26556
"111110000110000001110001100000000000",--26557
"111110000110100000000001100000000000",--26558
"011110000111000000000000000000000010",--26559
"101110000011111000000001100000000000",--26560
"000101000000000000000110011111000011",--26561
"111110000110011000000001100000000000",--26562
"001111000000000001110000000100000110",--26563
"111110001110001000110011100000000000",--26564
"001011000000000001110000000100000110",--26565
"001111000000000001110000000100000111",--26566
"111110001110001000110011100000000000",--26567
"001011000000000001110000000100000111",--26568
"001111000000000001110000000100001000",--26569
"111110001110001000110001100000000000",--26570
"001011000000000000110000000100001000",--26571
"001011000000000000000000000100011101",--26572
"001011000000000000000000000100011110",--26573
"001011000000000000000000000100011111",--26574
"001111000000000000110000000101100111",--26575
"001011000000000000110000000100010101",--26576
"001111000000000000110000000101101000",--26577
"001011000000000000110000000100010110",--26578
"001111000000000000110000000101101001",--26579
"001011000000000000110000000100010111",--26580
"101110000011111000000001100000000000",--26581
"001101111100000001011111111111111100",--26582
"001100001010000000010001100000000000",--26583
"001001111100000000101111111111111010",--26584
"001001111100000000011111111111111001",--26585
"101001000000000000100000000100000110",--26586
"101000000001111000000000100000000000",--26587
"101110000001111000000010000000000000",--26588
"001001111100000111111111111111111000",--26589
"101001111100010111100000000000001001",--26590
"000111000000000000000011010111001111",--26591
"101001111100000111100000000000001001",--26592
"001101111100000111111111111111111000",--26593
"001101111100000000011111111111111001",--26594
"001101111100000000111111111111111100",--26595
"001100000110000000010001000000000000",--26596
"001101000100000000100000000000000000",--26597
"001111000000000000110000000100011101",--26598
"001011000100000000110000000000000000",--26599
"001111000000000000110000000100011110",--26600
"001011000100000000110000000000000001",--26601
"001111000000000000110000000100011111",--26602
"001011000100000000110000000000000010",--26603
"001100000110000000010001000000000000",--26604
"001101000100000000100000000000000110",--26605
"001101111100000001001111111111111010",--26606
"001001000100000001000000000000000000",--26607
"001100000110000000010001000000000000",--26608
"001101000100000001010000000000000010",--26609
"001101001010000001100000000000000000",--26610
"010111001101000000000000000100101011",--26611
"001101000100000001100000000000000011",--26612
"001101001100000001110000000000000000",--26613
"001001111100000000101111111111111000",--26614
"001001111100000001101111111111110111",--26615
"001001111100000001011111111111110110",--26616
"010000001111000000000000000011111111",--26617
"001101000100000001110000000000000110",--26618
"001101001110000001110000000000000000",--26619
"001011000000000000000000000100100000",--26620
"001011000000000000000000000100100001",--26621
"001011000000000000000000000100100010",--26622
"001101000100000010000000000000000111",--26623
"001101000100000010010000000000000001",--26624
"001101001110000001110000000011111110",--26625
"001101010000000010000000000000000000",--26626
"001101010010000010010000000000000000",--26627
"001111010010000000110000000000000000",--26628
"001011000000000000110000000100010010",--26629
"001111010010000000110000000000000001",--26630
"001011000000000000110000000100010011",--26631
"001111010010000000110000000000000010",--26632
"001011000000000000110000000100010100",--26633
"001101000000000010100000000110101010",--26634
"101001010100010010100000000000000001",--26635
"001001111100000010011111111111110101",--26636
"001001111100000010001111111111110100",--26637
"001001111100000001111111111111110011",--26638
"010111010101000000000000000011010111",--26639
"001101010100000010110000000101101101",--26640
"001101010110000011000000000000001010",--26641
"001101010110000011010000000000000001",--26642
"001111010010000000110000000000000000",--26643
"001101010110000011100000000000000101",--26644
"001111011100000001000000000000000000",--26645
"111110000110010001000001100000000000",--26646
"001011011000000000110000000000000000",--26647
"001111010010000000110000000000000001",--26648
"001111011100000001000000000000000001",--26649
"111110000110010001000001100000000000",--26650
"001011011000000000110000000000000001",--26651
"001111010010000000110000000000000010",--26652
"001111011100000001000000000000000010",--26653
"111110000110010001000001100000000000",--26654
"001011011000000000110000000000000010",--26655
"011111011011000000100000000000001110",--26656
"001101010110000010110000000000000100",--26657
"001111011000000000110000000000000000",--26658
"001111011000000001000000000000000001",--26659
"001111011000000001010000000000000010",--26660
"001111010110000001100000000000000000",--26661
"111110001100001000110001100000000000",--26662
"001111010110000001100000000000000001",--26663
"111110001100001001000010000000000000",--26664
"111110000110000001000001100000000000",--26665
"001111010110000001000000000000000010",--26666
"111110001000001001010010000000000000",--26667
"111110000110000001000001100000000000",--26668
"001011011000000000110000000000000011",--26669
"000101000000000000000110100001010100",--26670
"010111011011000000100000000000100100",--26671
"001111011000000000110000000000000000",--26672
"001111011000000001000000000000000001",--26673
"001111011000000001010000000000000010",--26674
"111110000110001000110011000000000000",--26675
"001101010110000011100000000000000100",--26676
"001111011100000001110000000000000000",--26677
"111110001100001001110011000000000000",--26678
"111110001000001001000011100000000000",--26679
"001111011100000010000000000000000001",--26680
"111110001110001010000011100000000000",--26681
"111110001100000001110011000000000000",--26682
"111110001010001001010011100000000000",--26683
"001111011100000010000000000000000010",--26684
"111110001110001010000011100000000000",--26685
"111110001100000001110011000000000000",--26686
"001101010110000011100000000000000011",--26687
"011100011101000000000000000000000011",--26688
"101110001101111000000001100000000000",--26689
"011111011011000000110000000000010000",--26690
"000101000000000000000110100001010010",--26691
"111110001000001001010011100000000000",--26692
"001101010110000010110000000000001001",--26693
"001111010110000010000000000000000000",--26694
"111110001110001010000011100000000000",--26695
"111110001100000001110011000000000000",--26696
"111110001010001000110010100000000000",--26697
"001111010110000001110000000000000001",--26698
"111110001010001001110010100000000000",--26699
"111110001100000001010010100000000000",--26700
"111110000110001001000001100000000000",--26701
"001111010110000001000000000000000010",--26702
"111110000110001001000001100000000000",--26703
"111110001010000000110001100000000000",--26704
"011111011011000000110000000000000001",--26705
"111110000110010000010001100000000000",--26706
"001011011000000000110000000000000011",--26707
"101001010100010010100000000000000001",--26708
"010111010101000000000000000010010001",--26709
"001101010100000010110000000101101101",--26710
"001101010110000011000000000000001010",--26711
"001101010110000011010000000000000001",--26712
"001111010010000000110000000000000000",--26713
"001101010110000011100000000000000101",--26714
"001111011100000001000000000000000000",--26715
"111110000110010001000001100000000000",--26716
"001011011000000000110000000000000000",--26717
"001111010010000000110000000000000001",--26718
"001111011100000001000000000000000001",--26719
"111110000110010001000001100000000000",--26720
"001011011000000000110000000000000001",--26721
"001111010010000000110000000000000010",--26722
"001111011100000001000000000000000010",--26723
"111110000110010001000001100000000000",--26724
"001011011000000000110000000000000010",--26725
"011111011011000000100000000000001110",--26726
"001101010110000010110000000000000100",--26727
"001111011000000000110000000000000000",--26728
"001111011000000001000000000000000001",--26729
"001111011000000001010000000000000010",--26730
"001111010110000001100000000000000000",--26731
"111110001100001000110001100000000000",--26732
"001111010110000001100000000000000001",--26733
"111110001100001001000010000000000000",--26734
"111110000110000001000001100000000000",--26735
"001111010110000001000000000000000010",--26736
"111110001000001001010010000000000000",--26737
"111110000110000001000001100000000000",--26738
"001011011000000000110000000000000011",--26739
"000101000000000000000110100010011010",--26740
"010111011011000000100000000000100100",--26741
"001111011000000000110000000000000000",--26742
"001111011000000001000000000000000001",--26743
"001111011000000001010000000000000010",--26744
"111110000110001000110011000000000000",--26745
"001101010110000011100000000000000100",--26746
"001111011100000001110000000000000000",--26747
"111110001100001001110011000000000000",--26748
"111110001000001001000011100000000000",--26749
"001111011100000010000000000000000001",--26750
"111110001110001010000011100000000000",--26751
"111110001100000001110011000000000000",--26752
"111110001010001001010011100000000000",--26753
"001111011100000010000000000000000010",--26754
"111110001110001010000011100000000000",--26755
"111110001100000001110011000000000000",--26756
"001101010110000011100000000000000011",--26757
"011100011101000000000000000000000011",--26758
"101110001101111000000001100000000000",--26759
"011111011011000000110000000000010000",--26760
"000101000000000000000110100010011000",--26761
"111110001000001001010011100000000000",--26762
"001101010110000010110000000000001001",--26763
"001111010110000010000000000000000000",--26764
"111110001110001010000011100000000000",--26765
"111110001100000001110011000000000000",--26766
"111110001010001000110010100000000000",--26767
"001111010110000001110000000000000001",--26768
"111110001010001001110010100000000000",--26769
"111110001100000001010010100000000000",--26770
"111110000110001001000001100000000000",--26771
"001111010110000001000000000000000010",--26772
"111110000110001001000001100000000000",--26773
"111110001010000000110001100000000000",--26774
"011111011011000000110000000000000001",--26775
"111110000110010000010001100000000000",--26776
"001011011000000000110000000000000011",--26777
"101001010100010010100000000000000001",--26778
"010111010101000000000000000001001011",--26779
"001101010100000010110000000101101101",--26780
"001101010110000011000000000000001010",--26781
"001101010110000011010000000000000001",--26782
"001111010010000000110000000000000000",--26783
"001101010110000011100000000000000101",--26784
"001111011100000001000000000000000000",--26785
"111110000110010001000001100000000000",--26786
"001011011000000000110000000000000000",--26787
"001111010010000000110000000000000001",--26788
"001111011100000001000000000000000001",--26789
"111110000110010001000001100000000000",--26790
"001011011000000000110000000000000001",--26791
"001111010010000000110000000000000010",--26792
"001111011100000001000000000000000010",--26793
"111110000110010001000001100000000000",--26794
"001011011000000000110000000000000010",--26795
"011111011011000000100000000000001110",--26796
"001101010110000010110000000000000100",--26797
"001111011000000000110000000000000000",--26798
"001111011000000001000000000000000001",--26799
"001111011000000001010000000000000010",--26800
"001111010110000001100000000000000000",--26801
"111110001100001000110001100000000000",--26802
"001111010110000001100000000000000001",--26803
"111110001100001001000010000000000000",--26804
"111110000110000001000001100000000000",--26805
"001111010110000001000000000000000010",--26806
"111110001000001001010010000000000000",--26807
"111110000110000001000001100000000000",--26808
"001011011000000000110000000000000011",--26809
"000101000000000000000110100011100000",--26810
"010111011011000000100000000000100100",--26811
"001111011000000000110000000000000000",--26812
"001111011000000001000000000000000001",--26813
"001111011000000001010000000000000010",--26814
"111110000110001000110011000000000000",--26815
"001101010110000011100000000000000100",--26816
"001111011100000001110000000000000000",--26817
"111110001100001001110011000000000000",--26818
"111110001000001001000011100000000000",--26819
"001111011100000010000000000000000001",--26820
"111110001110001010000011100000000000",--26821
"111110001100000001110011000000000000",--26822
"111110001010001001010011100000000000",--26823
"001111011100000010000000000000000010",--26824
"111110001110001010000011100000000000",--26825
"111110001100000001110011000000000000",--26826
"001101010110000011100000000000000011",--26827
"011100011101000000000000000000000011",--26828
"101110001101111000000001100000000000",--26829
"011111011011000000110000000000010000",--26830
"000101000000000000000110100011011110",--26831
"111110001000001001010011100000000000",--26832
"001101010110000010110000000000001001",--26833
"001111010110000010000000000000000000",--26834
"111110001110001010000011100000000000",--26835
"111110001100000001110011000000000000",--26836
"111110001010001000110010100000000000",--26837
"001111010110000001110000000000000001",--26838
"111110001010001001110010100000000000",--26839
"111110001100000001010010100000000000",--26840
"111110000110001001000001100000000000",--26841
"001111010110000001000000000000000010",--26842
"111110000110001001000001100000000000",--26843
"111110001010000000110001100000000000",--26844
"011111011011000000110000000000000001",--26845
"111110000110010000010001100000000000",--26846
"001011011000000000110000000000000011",--26847
"101001010100010000100000000000000001",--26848
"101000010011111000000000100000000000",--26849
"001001111100000111111111111111110010",--26850
"101001111100010111100000000000001111",--26851
"000111000000000000000000011001101110",--26852
"101001111100000111100000000000001111",--26853
"001101111100000111111111111111110010",--26854
"101001000000000001000000000001110110",--26855
"001101111100000000011111111111110011",--26856
"001101111100000000101111111111110100",--26857
"001101111100000000111111111111110101",--26858
"001001111100000111111111111111110010",--26859
"101001111100010111100000000000001111",--26860
"000111000000000000000100000011011010",--26861
"101001111100000111100000000000001111",--26862
"001101111100000111111111111111110010",--26863
"001101111100000000011111111111111000",--26864
"001101000010000000100000000000000101",--26865
"001101000100000000100000000000000000",--26866
"001111000000000000110000000100100000",--26867
"001011000100000000110000000000000000",--26868
"001111000000000000110000000100100001",--26869
"001011000100000000110000000000000001",--26870
"001111000000000000110000000100100010",--26871
"001011000100000000110000000000000010",--26872
"001101111100000000011111111111110110",--26873
"001101000010000000010000000000000001",--26874
"010111000011000000000000000000100011",--26875
"001101111100000000011111111111110111",--26876
"001101000010000000010000000000000001",--26877
"010000000011000000000000000000011001",--26878
"001101111100000000011111111111111000",--26879
"001101000010000000100000000000000110",--26880
"001101000100000000100000000000000000",--26881
"001011000000000000000000000100100000",--26882
"001011000000000000000000000100100001",--26883
"001011000000000000000000000100100010",--26884
"001101000010000000110000000000000111",--26885
"001101000010000001000000000000000001",--26886
"001101000100000000010000000011111110",--26887
"001101000110000000100000000000000001",--26888
"001101001000000000110000000000000001",--26889
"001001111100000111111111111111110101",--26890
"101001111100010111100000000000001100",--26891
"000111000000000000000100101110010000",--26892
"101001111100000111100000000000001100",--26893
"001101111100000111111111111111110101",--26894
"001101111100000000011111111111111000",--26895
"001101000010000000100000000000000101",--26896
"001101000100000000100000000000000001",--26897
"001111000000000000110000000100100000",--26898
"001011000100000000110000000000000000",--26899
"001111000000000000110000000100100001",--26900
"001011000100000000110000000000000001",--26901
"001111000000000000110000000100100010",--26902
"001011000100000000110000000000000010",--26903
"101001000000000000100000000000000010",--26904
"001101111100000000011111111111111000",--26905
"001001111100000111111111111111110101",--26906
"101001111100010111100000000000001100",--26907
"000111000000000000000110001000010000",--26908
"101001111100000111100000000000001100",--26909
"001101111100000111111111111111110101",--26910
"001101111100000000011111111111111001",--26911
"101001000010010000100000000000000001",--26912
"001101111100000000011111111111111010",--26913
"101001000010000000010000000000000001",--26914
"011011000011000001010000000000000010",--26915
"101000000011111000000001100000000000",--26916
"000101000000000000000110100100100111",--26917
"101001000010010000110000000000000101",--26918
"001111111100000000111111111111111110",--26919
"001111111100000001001111111111111111",--26920
"001111111100000001010000000000000000",--26921
"001101111100000000011111111111111100",--26922
"010111000100000000001111100000000000",--26923
"000101000000000000000110010100111010",--26924
"001101000000000001100000000100011011",--26925
"010100001100000000011111100000000000",--26926
"001100001000000000010011000000000000",--26927
"001101001100000001100000000000000000",--26928
"001111001100000000110000000000000000",--26929
"001011000000000000110000000100011101",--26930
"001111001100000000110000000000000001",--26931
"001011000000000000110000000100011110",--26932
"001111001100000000110000000000000010",--26933
"001011000000000000110000000100011111",--26934
"001101000000000001100000000100011100",--26935
"101001000100000001110000000000000001",--26936
"010100001101000001110000000000001101",--26937
"010100000101000000000000000000001010",--26938
"001101000000000001100000000100011011",--26939
"101001000010000001110000000000000001",--26940
"010100001101000001110000000000000101",--26941
"010100000011000000000000000000000010",--26942
"101001000000000001100000000000000001",--26943
"000101000000000000000110100101001000",--26944
"101000000001111000000011000000000000",--26945
"000101000000000000000110100101001000",--26946
"101000000001111000000011000000000000",--26947
"000101000000000000000110100101001000",--26948
"101000000001111000000011000000000000",--26949
"000101000000000000000110100101001000",--26950
"101000000001111000000011000000000000",--26951
"001001111100000001010000000000000000",--26952
"001001111100000001001111111111111111",--26953
"001001111100000000111111111111111110",--26954
"001001111100000000101111111111111101",--26955
"001001111100000000011111111111111100",--26956
"011100001101000000000000000010100111",--26957
"001100001000000000010011000000000000",--26958
"001101001100000001110000000000000010",--26959
"001101001110000010000000000000000000",--26960
"010111010001000000000000000101101001",--26961
"001101001100000010000000000000000011",--26962
"001101010000000010010000000000000000",--26963
"001001111100000001101111111111111011",--26964
"001001111100000010001111111111111010",--26965
"001001111100000001111111111111111001",--26966
"010000010011000000000000000001011000",--26967
"001101001100000010010000000000000101",--26968
"001101001100000010100000000000000111",--26969
"001101001100000010110000000000000001",--26970
"001101001100000011000000000000000100",--26971
"001101010010000010010000000000000000",--26972
"001111010010000000110000000000000000",--26973
"001011000000000000110000000100100000",--26974
"001111010010000000110000000000000001",--26975
"001011000000000000110000000100100001",--26976
"001111010010000000110000000000000010",--26977
"001011000000000000110000000100100010",--26978
"001101001100000010010000000000000110",--26979
"001101010010000010010000000000000000",--26980
"001101010100000010100000000000000000",--26981
"001101010110000010110000000000000000",--26982
"001001111100000011001111111111111000",--26983
"001001111100000010111111111111110111",--26984
"001001111100000010101111111111110110",--26985
"001001111100000010011111111111110101",--26986
"010000010011000000000000000000001000",--26987
"001101000000000000010000000011111110",--26988
"101000010111111000000001100000000000",--26989
"101000010101111000000001000000000000",--26990
"001001111100000111111111111111110100",--26991
"101001111100010111100000000000001101",--26992
"000111000000000000000100101110010000",--26993
"101001111100000111100000000000001101",--26994
"001101111100000111111111111111110100",--26995
"001101111100000000011111111111110101",--26996
"010011000011000000010000000000001000",--26997
"001101000000000000010000000011111111",--26998
"001101111100000000101111111111110110",--26999
"001101111100000000111111111111110111",--27000
"001001111100000111111111111111110100",--27001
"101001111100010111100000000000001101",--27002
"000111000000000000000100101110010000",--27003
"101001111100000111100000000000001101",--27004
"001101111100000111111111111111110100",--27005
"001101111100000000011111111111110101",--27006
"010011000011000000100000000000001000",--27007
"001101000000000000010000000100000000",--27008
"001101111100000000101111111111110110",--27009
"001101111100000000111111111111110111",--27010
"001001111100000111111111111111110100",--27011
"101001111100010111100000000000001101",--27012
"000111000000000000000100101110010000",--27013
"101001111100000111100000000000001101",--27014
"001101111100000111111111111111110100",--27015
"001101111100000000011111111111110101",--27016
"010011000011000000110000000000001000",--27017
"001101000000000000010000000100000001",--27018
"001101111100000000101111111111110110",--27019
"001101111100000000111111111111110111",--27020
"001001111100000111111111111111110100",--27021
"101001111100010111100000000000001101",--27022
"000111000000000000000100101110010000",--27023
"101001111100000111100000000000001101",--27024
"001101111100000111111111111111110100",--27025
"001101111100000000011111111111110101",--27026
"010011000011000001000000000000001000",--27027
"001101000000000000010000000100000010",--27028
"001101111100000000101111111111110110",--27029
"001101111100000000111111111111110111",--27030
"001001111100000111111111111111110100",--27031
"101001111100010111100000000000001101",--27032
"000111000000000000000100101110010000",--27033
"101001111100000111100000000000001101",--27034
"001101111100000111111111111111110100",--27035
"001101111100000000011111111111111000",--27036
"001101000010000000010000000000000000",--27037
"001111000000000000110000000100011101",--27038
"001111000010000001000000000000000000",--27039
"001111000000000001010000000100100000",--27040
"111110001000001001010010000000000000",--27041
"111110000110000001000001100000000000",--27042
"001011000000000000110000000100011101",--27043
"001111000000000000110000000100011110",--27044
"001111000010000001000000000000000001",--27045
"001111000000000001010000000100100001",--27046
"111110001000001001010010000000000000",--27047
"111110000110000001000001100000000000",--27048
"001011000000000000110000000100011110",--27049
"001111000000000000110000000100011111",--27050
"001111000010000001000000000000000010",--27051
"001111000000000001010000000100100010",--27052
"111110001000001001010010000000000000",--27053
"111110000110000001000001100000000000",--27054
"001011000000000000110000000100011111",--27055
"001101111100000000011111111111111001",--27056
"001101000010000000100000000000000001",--27057
"010111000101000000000000000100001000",--27058
"001101111100000000101111111111111010",--27059
"001101000100000000110000000000000001",--27060
"010000000111000000000000000000101010",--27061
"001101111100000000111111111111111011",--27062
"001101000110000001000000000000000101",--27063
"001101000110000001010000000000000111",--27064
"001101000110000001100000000000000001",--27065
"001101000110000001110000000000000100",--27066
"001101001000000001000000000000000001",--27067
"001111001000000000110000000000000000",--27068
"001011000000000000110000000100100000",--27069
"001111001000000000110000000000000001",--27070
"001011000000000000110000000100100001",--27071
"001111001000000000110000000000000010",--27072
"001011000000000000110000000100100010",--27073
"001101000110000001000000000000000110",--27074
"001101001000000000010000000000000000",--27075
"001101001010000000100000000000000001",--27076
"001101001100000000110000000000000001",--27077
"001001111100000001111111111111111000",--27078
"001001111100000111111111111111110111",--27079
"101001111100010111100000000000001010",--27080
"000111000000000000000101000111001101",--27081
"101001111100000111100000000000001010",--27082
"001101111100000111111111111111110111",--27083
"001101111100000000011111111111111000",--27084
"001101000010000000010000000000000001",--27085
"001111000000000000110000000100011101",--27086
"001111000010000001000000000000000000",--27087
"001111000000000001010000000100100000",--27088
"111110001000001001010010000000000000",--27089
"111110000110000001000001100000000000",--27090
"001011000000000000110000000100011101",--27091
"001111000000000000110000000100011110",--27092
"001111000010000001000000000000000001",--27093
"001111000000000001010000000100100001",--27094
"111110001000001001010010000000000000",--27095
"111110000110000001000001100000000000",--27096
"001011000000000000110000000100011110",--27097
"001111000000000000110000000100011111",--27098
"001111000010000001000000000000000010",--27099
"001111000000000001010000000100100010",--27100
"111110001000001001010010000000000000",--27101
"111110000110000001000001100000000000",--27102
"001011000000000000110000000100011111",--27103
"101001000000000000100000000000000010",--27104
"001101111100000000011111111111111001",--27105
"001101000010000000010000000000000010",--27106
"010111000011000000000000000011010111",--27107
"001101111100000000011111111111111010",--27108
"001101000010000000010000000000000010",--27109
"010000000011000000000000000000000110",--27110
"001101111100000000011111111111111011",--27111
"001001111100000111111111111111111000",--27112
"101001111100010111100000000000001001",--27113
"000111000000000000000101011001110000",--27114
"101001111100000111100000000000001001",--27115
"001101111100000111111111111111111000",--27116
"101001000000000000100000000000000011",--27117
"001101111100000000011111111111111011",--27118
"001001111100000111111111111111111000",--27119
"101001111100010111100000000000001001",--27120
"000111000000000000000101101010010000",--27121
"101001111100000111100000000000001001",--27122
"001101111100000111111111111111111000",--27123
"000101000000000000000110101010111011",--27124
"001100001000000000010011000000000000",--27125
"001101001100000001110000000000000010",--27126
"001101001110000001110000000000000000",--27127
"010111001111000000000000000011000010",--27128
"001100001000000000010011100000000000",--27129
"001101001110000001110000000000000010",--27130
"001101001110000001110000000000000000",--27131
"001100000110000000010100000000000000",--27132
"001101010000000010000000000000000010",--27133
"001101010000000010000000000000000000",--27134
"011100010001000001110000000000001110",--27135
"001100001010000000010100000000000000",--27136
"001101010000000010000000000000000010",--27137
"001101010000000010000000000000000000",--27138
"011100010001000001110000000000001010",--27139
"101001000010010010000000000000000001",--27140
"001100001000000010000100000000000000",--27141
"001101010000000010000000000000000010",--27142
"001101010000000010000000000000000000",--27143
"011100010001000001110000000000000101",--27144
"101001000010000010000000000000000001",--27145
"001100001000000010000100000000000000",--27146
"001101010000000010000000000000000010",--27147
"001101010000000010000000000000000000",--27148
"010000010001000001110000000001001000",--27149
"001100001000000000010011000000000000",--27150
"001101001100000001110000000000000010",--27151
"001101001110000010000000000000000000",--27152
"010111010001000000000000000010101001",--27153
"001101001100000010000000000000000011",--27154
"001101010000000010010000000000000000",--27155
"001001111100000001101111111111111011",--27156
"001001111100000010001111111111111010",--27157
"001001111100000001111111111111111001",--27158
"010000010011000000000000000000101001",--27159
"001101001100000010010000000000000101",--27160
"001101001100000010100000000000000111",--27161
"001101001100000010110000000000000001",--27162
"001101001100000011000000000000000100",--27163
"001101010010000010010000000000000000",--27164
"001111010010000000110000000000000000",--27165
"001011000000000000110000000100100000",--27166
"001111010010000000110000000000000001",--27167
"001011000000000000110000000100100001",--27168
"001111010010000000110000000000000010",--27169
"001011000000000000110000000100100010",--27170
"001101001100000010010000000000000110",--27171
"001101010010000000010000000000000000",--27172
"001101010100000000100000000000000000",--27173
"001101010110000000110000000000000000",--27174
"001001111100000011001111111111111000",--27175
"001001111100000111111111111111110111",--27176
"101001111100010111100000000000001010",--27177
"000111000000000000000101000111001101",--27178
"101001111100000111100000000000001010",--27179
"001101111100000111111111111111110111",--27180
"001101111100000000011111111111111000",--27181
"001101000010000000010000000000000000",--27182
"001111000000000000110000000100011101",--27183
"001111000010000001000000000000000000",--27184
"001111000000000001010000000100100000",--27185
"111110001000001001010010000000000000",--27186
"111110000110000001000001100000000000",--27187
"001011000000000000110000000100011101",--27188
"001111000000000000110000000100011110",--27189
"001111000010000001000000000000000001",--27190
"001111000000000001010000000100100001",--27191
"111110001000001001010010000000000000",--27192
"111110000110000001000001100000000000",--27193
"001011000000000000110000000100011110",--27194
"001111000000000000110000000100011111",--27195
"001111000010000001000000000000000010",--27196
"001111000000000001010000000100100010",--27197
"111110001000001001010010000000000000",--27198
"111110000110000001000001100000000000",--27199
"001011000000000000110000000100011111",--27200
"101001000000000000100000000000000001",--27201
"001101111100000000011111111111111001",--27202
"001101000010000000010000000000000001",--27203
"010111000011000000000000000001110110",--27204
"001101111100000000011111111111111010",--27205
"001101000010000000010000000000000001",--27206
"010000000011000000000000000000000110",--27207
"001101111100000000011111111111111011",--27208
"001001111100000111111111111111111000",--27209
"101001111100010111100000000000001001",--27210
"000111000000000000000101011001110000",--27211
"101001111100000111100000000000001001",--27212
"001101111100000111111111111111111000",--27213
"101001000000000000100000000000000010",--27214
"001101111100000000011111111111111011",--27215
"001001111100000111111111111111111000",--27216
"101001111100010111100000000000001001",--27217
"000111000000000000000101101010010000",--27218
"101001111100000111100000000000001001",--27219
"001101111100000111111111111111111000",--27220
"000101000000000000000110101010111011",--27221
"001101001100000001100000000000000011",--27222
"001101001100000001100000000000000000",--27223
"010000001101000000000000000001011100",--27224
"001100000110000000010011000000000000",--27225
"001101001100000001100000000000000101",--27226
"101001000010010001110000000000000001",--27227
"001100001000000001110011100000000000",--27228
"001101001110000001110000000000000101",--27229
"001100001000000000010100000000000000",--27230
"001101010000000010000000000000000101",--27231
"101001000010000010010000000000000001",--27232
"001100001000000010010100100000000000",--27233
"001101010010000010010000000000000101",--27234
"001100001010000000010101000000000000",--27235
"001101010100000010100000000000000101",--27236
"001101001100000001100000000000000000",--27237
"001111001100000000110000000000000000",--27238
"001011000000000000110000000100100000",--27239
"001111001100000000110000000000000001",--27240
"001011000000000000110000000100100001",--27241
"001111001100000000110000000000000010",--27242
"001011000000000000110000000100100010",--27243
"001101001110000001100000000000000000",--27244
"001111000000000000110000000100100000",--27245
"001111001100000001000000000000000000",--27246
"111110000110000001000001100000000000",--27247
"001011000000000000110000000100100000",--27248
"001111000000000000110000000100100001",--27249
"001111001100000001000000000000000001",--27250
"111110000110000001000001100000000000",--27251
"001011000000000000110000000100100001",--27252
"001111000000000000110000000100100010",--27253
"001111001100000001000000000000000010",--27254
"111110000110000001000001100000000000",--27255
"001011000000000000110000000100100010",--27256
"001101010000000001100000000000000000",--27257
"001111000000000000110000000100100000",--27258
"001111001100000001000000000000000000",--27259
"111110000110000001000001100000000000",--27260
"001011000000000000110000000100100000",--27261
"001111000000000000110000000100100001",--27262
"001111001100000001000000000000000001",--27263
"111110000110000001000001100000000000",--27264
"001011000000000000110000000100100001",--27265
"001111000000000000110000000100100010",--27266
"001111001100000001000000000000000010",--27267
"111110000110000001000001100000000000",--27268
"001011000000000000110000000100100010",--27269
"001101010010000001100000000000000000",--27270
"001111000000000000110000000100100000",--27271
"001111001100000001000000000000000000",--27272
"111110000110000001000001100000000000",--27273
"001011000000000000110000000100100000",--27274
"001111000000000000110000000100100001",--27275
"001111001100000001000000000000000001",--27276
"111110000110000001000001100000000000",--27277
"001011000000000000110000000100100001",--27278
"001111000000000000110000000100100010",--27279
"001111001100000001000000000000000010",--27280
"111110000110000001000001100000000000",--27281
"001011000000000000110000000100100010",--27282
"001101010100000001100000000000000000",--27283
"001111000000000000110000000100100000",--27284
"001111001100000001000000000000000000",--27285
"111110000110000001000001100000000000",--27286
"001011000000000000110000000100100000",--27287
"001111000000000000110000000100100001",--27288
"001111001100000001000000000000000001",--27289
"111110000110000001000001100000000000",--27290
"001011000000000000110000000100100001",--27291
"001111000000000000110000000100100010",--27292
"001111001100000001000000000000000010",--27293
"111110000110000001000001100000000000",--27294
"001011000000000000110000000100100010",--27295
"001100001000000000010011000000000000",--27296
"001101001100000001100000000000000100",--27297
"001101001100000001100000000000000000",--27298
"001111000000000000110000000100011101",--27299
"001111001100000001000000000000000000",--27300
"001111000000000001010000000100100000",--27301
"111110001000001001010010000000000000",--27302
"111110000110000001000001100000000000",--27303
"001011000000000000110000000100011101",--27304
"001111000000000000110000000100011110",--27305
"001111001100000001000000000000000001",--27306
"001111000000000001010000000100100001",--27307
"111110001000001001010010000000000000",--27308
"111110000110000001000001100000000000",--27309
"001011000000000000110000000100011110",--27310
"001111000000000000110000000100011111",--27311
"001111001100000001000000000000000010",--27312
"001111000000000001010000000100100010",--27313
"111110001000001001010010000000000000",--27314
"111110000110000001000001100000000000",--27315
"001011000000000000110000000100011111",--27316
"101001000000000001100000000000000001",--27317
"001001111100000111111111111111111011",--27318
"101001111100010111100000000000000110",--27319
"000111000000000000000110000000010100",--27320
"101001111100000111100000000000000110",--27321
"001101111100000111111111111111111011",--27322
"001111000000000000110000000100011101",--27323
"101100000111101000000000100000000000",--27324
"010111000011111111110000000000000010",--27325
"101001000000000000010000000011111111",--27326
"000101000000000000000110101011000010",--27327
"011000000011000000000000000000000001",--27328
"101000000001111000000000100000000000",--27329
"000000000010000000000000000000000000",--27330
"001111000000000000110000000100011110",--27331
"101100000111101000000000100000000000",--27332
"010111000011111111110000000000000010",--27333
"101001000000000000010000000011111111",--27334
"000101000000000000000110101011001010",--27335
"011000000011000000000000000000000001",--27336
"101000000001111000000000100000000000",--27337
"000000000010000000000000000000000000",--27338
"001111000000000000110000000100011111",--27339
"101100000111101000000000100000000000",--27340
"010111000011111111110000000000000010",--27341
"101001000000000000010000000011111111",--27342
"000101000000000000000110101011010010",--27343
"011000000011000000000000000000000001",--27344
"101000000001111000000000100000000000",--27345
"000000000010000000000000000000000000",--27346
"001101111100000000011111111111111100",--27347
"101001000010000000010000000000000001",--27348
"001101111100000000101111111111111101",--27349
"001101111100000000111111111111111110",--27350
"001101111100000001001111111111111111",--27351
"001101111100000001010000000000000000",--27352
"000101000000000000000110100100101101",--27353
"001101000000000001100000000100011100",--27354
"010100001100000000011111100000000000",--27355
"101001001100010001100000000000000001",--27356
"001001111100000001010000000000000000",--27357
"001001111100000001001111111111111111",--27358
"001001111100000000111111111111111110",--27359
"001001111100000000101111111111111101",--27360
"001001111100000000011111111111111100",--27361
"010100001101000000010000000000011111",--27362
"101001000010000001100000000000000001",--27363
"001111000000000000110000000100011000",--27364
"001101000000000001110000000100011010",--27365
"101000001100010001110011000000000000",--27366
"101010001101101000000010000000000000",--27367
"111110000110001001000001100000000000",--27368
"001111000000000001000000000100001100",--27369
"111110000110001001000010000000000000",--27370
"001111000000000001010000000100001001",--27371
"111110001000000001010010000000000000",--27372
"001111000000000001010000000100001101",--27373
"111110000110001001010010100000000000",--27374
"001111000000000001100000000100001010",--27375
"111110001010000001100010100000000000",--27376
"001111000000000001100000000100001110",--27377
"111110000110001001100001100000000000",--27378
"001111000000000001100000000100001011",--27379
"111110000110000001100001100000000000",--27380
"001101000000000001100000000100011011",--27381
"101001001100010000100000000000000001",--27382
"101000001011111000000001100000000000",--27383
"101000001001111000000000100000000000",--27384
"101110001011111000001111100000000000",--27385
"101110000111111000000010100000000000",--27386
"101110001001111000000001100000000000",--27387
"101110111111111000000010000000000000",--27388
"001001111100000111111111111111111011",--27389
"101001111100010111100000000000000110",--27390
"000111000000000000000110010100111001",--27391
"101001111100000111100000000000000110",--27392
"001101111100000111111111111111111011",--27393
"101000000001111000000000100000000000",--27394
"001101111100000000101111111111111100",--27395
"001101111100000000111111111111111101",--27396
"001101111100000001001111111111111110",--27397
"001101111100000001011111111111111111",--27398
"001001111100000111111111111111111011",--27399
"101001111100010111100000000000000110",--27400
"000111000000000000000110100100101101",--27401
"101001111100000111100000000000000110",--27402
"001101111100000111111111111111111011",--27403
"001101111100000000011111111111111100",--27404
"101001000010000000010000000000000001",--27405
"001101111100000000100000000000000000",--27406
"101001000100000000100000000000000010",--27407
"011011000101000001010000000000000010",--27408
"101000000101111000000010100000000000",--27409
"000101000000000000000110101100010100",--27410
"101001000100010001010000000000000101",--27411
"001101111100000000101111111111111110",--27412
"001101111100000000111111111111111111",--27413
"001101111100000001001111111111111101",--27414
"000101000000000000000110101011011010",--27415
"101110000001111000000001100000000000",--27416
"001001111100000000010000000000000000",--27417
"001001111100000000101111111111111111",--27418
"101001000000000000010000000000000011",--27419
"001001111100000111111111111111111110",--27420
"000111000000000000000111010110110001",--27421
"001101111100000111111111111111111110",--27422
"101110000001111000000001100000000000",--27423
"001001111100000000011111111111111110",--27424
"101001000000000000010000000000000011",--27425
"001001111100000111111111111111111101",--27426
"000111000000000000000111010110110001",--27427
"101000000011111000000001000000000000",--27428
"101001000000000000010000000000000101",--27429
"000111000000000000000111010110101010",--27430
"001101111100000111111111111111111101",--27431
"101110000001111000000001100000000000",--27432
"001001111100000000011111111111111101",--27433
"101001000000000000010000000000000011",--27434
"001001111100000111111111111111111100",--27435
"000111000000000000000111010110110001",--27436
"001101111100000000101111111111111101",--27437
"001001000100000000010000000000000001",--27438
"101001000000000000010000000000000011",--27439
"101110000001111000000001100000000000",--27440
"000111000000000000000111010110110001",--27441
"001101111100000000101111111111111101",--27442
"001001000100000000010000000000000010",--27443
"101001000000000000010000000000000011",--27444
"101110000001111000000001100000000000",--27445
"000111000000000000000111010110110001",--27446
"001101111100000000101111111111111101",--27447
"001001000100000000010000000000000011",--27448
"101001000000000000010000000000000011",--27449
"101110000001111000000001100000000000",--27450
"000111000000000000000111010110110001",--27451
"001101111100000000101111111111111101",--27452
"001001000100000000010000000000000100",--27453
"101001000000000000010000000000000101",--27454
"101000000001111000000001000000000000",--27455
"000111000000000000000111010110101010",--27456
"001101111100000111111111111111111100",--27457
"001001111100000000011111111111111100",--27458
"101001000000000000010000000000000101",--27459
"101000000001111000000001000000000000",--27460
"001001111100000111111111111111111011",--27461
"000111000000000000000111010110101010",--27462
"001101111100000111111111111111111011",--27463
"101110000001111000000001100000000000",--27464
"001001111100000000011111111111111011",--27465
"101001000000000000010000000000000011",--27466
"001001111100000111111111111111111010",--27467
"000111000000000000000111010110110001",--27468
"101000000011111000000001000000000000",--27469
"101001000000000000010000000000000101",--27470
"000111000000000000000111010110101010",--27471
"001101111100000111111111111111111010",--27472
"101110000001111000000001100000000000",--27473
"001001111100000000011111111111111010",--27474
"101001000000000000010000000000000011",--27475
"001001111100000111111111111111111001",--27476
"000111000000000000000111010110110001",--27477
"001101111100000000101111111111111010",--27478
"001001000100000000010000000000000001",--27479
"101001000000000000010000000000000011",--27480
"101110000001111000000001100000000000",--27481
"000111000000000000000111010110110001",--27482
"001101111100000000101111111111111010",--27483
"001001000100000000010000000000000010",--27484
"101001000000000000010000000000000011",--27485
"101110000001111000000001100000000000",--27486
"000111000000000000000111010110110001",--27487
"001101111100000000101111111111111010",--27488
"001001000100000000010000000000000011",--27489
"101001000000000000010000000000000011",--27490
"101110000001111000000001100000000000",--27491
"000111000000000000000111010110110001",--27492
"001101111100000000101111111111111010",--27493
"001001000100000000010000000000000100",--27494
"101001000000000000010000000000000011",--27495
"101110000001111000000001100000000000",--27496
"000111000000000000000111010110110001",--27497
"101000000011111000000001000000000000",--27498
"101001000000000000010000000000000101",--27499
"000111000000000000000111010110101010",--27500
"001101111100000111111111111111111001",--27501
"101110000001111000000001100000000000",--27502
"001001111100000000011111111111111001",--27503
"101001000000000000010000000000000011",--27504
"001001111100000111111111111111111000",--27505
"000111000000000000000111010110110001",--27506
"001101111100000000101111111111111001",--27507
"001001000100000000010000000000000001",--27508
"101001000000000000010000000000000011",--27509
"101110000001111000000001100000000000",--27510
"000111000000000000000111010110110001",--27511
"001101111100000000101111111111111001",--27512
"001001000100000000010000000000000010",--27513
"101001000000000000010000000000000011",--27514
"101110000001111000000001100000000000",--27515
"000111000000000000000111010110110001",--27516
"001101111100000000101111111111111001",--27517
"001001000100000000010000000000000011",--27518
"101001000000000000010000000000000011",--27519
"101110000001111000000001100000000000",--27520
"000111000000000000000111010110110001",--27521
"001101111100000000101111111111111001",--27522
"001001000100000000010000000000000100",--27523
"101001000000000000010000000000000001",--27524
"101000000001111000000001000000000000",--27525
"000111000000000000000111010110101010",--27526
"001101111100000111111111111111111000",--27527
"101110000001111000000001100000000000",--27528
"001001111100000000011111111111111000",--27529
"101001000000000000010000000000000011",--27530
"001001111100000111111111111111110111",--27531
"000111000000000000000111010110110001",--27532
"101000000011111000000001000000000000",--27533
"101001000000000000010000000000000101",--27534
"000111000000000000000111010110101010",--27535
"001101111100000111111111111111110111",--27536
"101110000001111000000001100000000000",--27537
"001001111100000000011111111111110111",--27538
"101001000000000000010000000000000011",--27539
"001001111100000111111111111111110110",--27540
"000111000000000000000111010110110001",--27541
"001101111100000000101111111111110111",--27542
"001001000100000000010000000000000001",--27543
"101001000000000000010000000000000011",--27544
"101110000001111000000001100000000000",--27545
"000111000000000000000111010110110001",--27546
"001101111100000000101111111111110111",--27547
"001001000100000000010000000000000010",--27548
"101001000000000000010000000000000011",--27549
"101110000001111000000001100000000000",--27550
"000111000000000000000111010110110001",--27551
"001101111100000000101111111111110111",--27552
"001001000100000000010000000000000011",--27553
"101001000000000000010000000000000011",--27554
"101110000001111000000001100000000000",--27555
"000111000000000000000111010110110001",--27556
"001101111100000111111111111111110110",--27557
"001101111100000000101111111111110111",--27558
"001001000100000000010000000000000100",--27559
"101000111011111000000000100000000000",--27560
"101001111010000111010000000000001000",--27561
"001001000010000000100000000000000111",--27562
"001101111100000000101111111111111000",--27563
"001001000010000000100000000000000110",--27564
"001101111100000000101111111111111001",--27565
"001001000010000000100000000000000101",--27566
"001101111100000000101111111111111010",--27567
"001001000010000000100000000000000100",--27568
"001101111100000000101111111111111011",--27569
"001001000010000000100000000000000011",--27570
"001101111100000000101111111111111100",--27571
"001001000010000000100000000000000010",--27572
"001101111100000000101111111111111101",--27573
"001001000010000000100000000000000001",--27574
"001101111100000000101111111111111110",--27575
"001001000010000000100000000000000000",--27576
"001101111100000000101111111111111111",--27577
"001101111100000001000000000000000000",--27578
"001000001000000000100000100000000000",--27579
"101001000100010000100000000000000001",--27580
"101000001001111000000000100000000000",--27581
"010111000100000000001111100000000000",--27582
"000101000000000000000110101100011000",--27583
"001101000000000000010000000100011011",--27584
"101110000001111000000001100000000000",--27585
"001001111100000000010000000000000000",--27586
"101001000000000000010000000000000011",--27587
"001001111100000111111111111111111111",--27588
"000111000000000000000111010110110001",--27589
"001101111100000111111111111111111111",--27590
"101110000001111000000001100000000000",--27591
"001001111100000000011111111111111111",--27592
"101001000000000000010000000000000011",--27593
"001001111100000111111111111111111110",--27594
"000111000000000000000111010110110001",--27595
"101000000011111000000001000000000000",--27596
"101001000000000000010000000000000101",--27597
"000111000000000000000111010110101010",--27598
"001101111100000111111111111111111110",--27599
"101110000001111000000001100000000000",--27600
"001001111100000000011111111111111110",--27601
"101001000000000000010000000000000011",--27602
"001001111100000111111111111111111101",--27603
"000111000000000000000111010110110001",--27604
"001101111100000000101111111111111110",--27605
"001001000100000000010000000000000001",--27606
"101001000000000000010000000000000011",--27607
"101110000001111000000001100000000000",--27608
"000111000000000000000111010110110001",--27609
"001101111100000000101111111111111110",--27610
"001001000100000000010000000000000010",--27611
"101001000000000000010000000000000011",--27612
"101110000001111000000001100000000000",--27613
"000111000000000000000111010110110001",--27614
"001101111100000000101111111111111110",--27615
"001001000100000000010000000000000011",--27616
"101001000000000000010000000000000011",--27617
"101110000001111000000001100000000000",--27618
"000111000000000000000111010110110001",--27619
"001101111100000000101111111111111110",--27620
"001001000100000000010000000000000100",--27621
"101001000000000000010000000000000101",--27622
"101000000001111000000001000000000000",--27623
"000111000000000000000111010110101010",--27624
"001101111100000111111111111111111101",--27625
"001001111100000000011111111111111101",--27626
"101001000000000000010000000000000101",--27627
"101000000001111000000001000000000000",--27628
"001001111100000111111111111111111100",--27629
"000111000000000000000111010110101010",--27630
"001101111100000111111111111111111100",--27631
"101110000001111000000001100000000000",--27632
"001001111100000000011111111111111100",--27633
"101001000000000000010000000000000011",--27634
"001001111100000111111111111111111011",--27635
"000111000000000000000111010110110001",--27636
"101000000011111000000001000000000000",--27637
"101001000000000000010000000000000101",--27638
"000111000000000000000111010110101010",--27639
"001101111100000111111111111111111011",--27640
"101110000001111000000001100000000000",--27641
"001001111100000000011111111111111011",--27642
"101001000000000000010000000000000011",--27643
"001001111100000111111111111111111010",--27644
"000111000000000000000111010110110001",--27645
"001101111100000000101111111111111011",--27646
"001001000100000000010000000000000001",--27647
"101001000000000000010000000000000011",--27648
"101110000001111000000001100000000000",--27649
"000111000000000000000111010110110001",--27650
"001101111100000000101111111111111011",--27651
"001001000100000000010000000000000010",--27652
"101001000000000000010000000000000011",--27653
"101110000001111000000001100000000000",--27654
"000111000000000000000111010110110001",--27655
"001101111100000000101111111111111011",--27656
"001001000100000000010000000000000011",--27657
"101001000000000000010000000000000011",--27658
"101110000001111000000001100000000000",--27659
"000111000000000000000111010110110001",--27660
"001101111100000000101111111111111011",--27661
"001001000100000000010000000000000100",--27662
"101001000000000000010000000000000011",--27663
"101110000001111000000001100000000000",--27664
"000111000000000000000111010110110001",--27665
"101000000011111000000001000000000000",--27666
"101001000000000000010000000000000101",--27667
"000111000000000000000111010110101010",--27668
"001101111100000111111111111111111010",--27669
"101110000001111000000001100000000000",--27670
"001001111100000000011111111111111010",--27671
"101001000000000000010000000000000011",--27672
"001001111100000111111111111111111001",--27673
"000111000000000000000111010110110001",--27674
"001101111100000000101111111111111010",--27675
"001001000100000000010000000000000001",--27676
"101001000000000000010000000000000011",--27677
"101110000001111000000001100000000000",--27678
"000111000000000000000111010110110001",--27679
"001101111100000000101111111111111010",--27680
"001001000100000000010000000000000010",--27681
"101001000000000000010000000000000011",--27682
"101110000001111000000001100000000000",--27683
"000111000000000000000111010110110001",--27684
"001101111100000000101111111111111010",--27685
"001001000100000000010000000000000011",--27686
"101001000000000000010000000000000011",--27687
"101110000001111000000001100000000000",--27688
"000111000000000000000111010110110001",--27689
"001101111100000000101111111111111010",--27690
"001001000100000000010000000000000100",--27691
"101001000000000000010000000000000001",--27692
"101000000001111000000001000000000000",--27693
"000111000000000000000111010110101010",--27694
"001101111100000111111111111111111001",--27695
"101110000001111000000001100000000000",--27696
"001001111100000000011111111111111001",--27697
"101001000000000000010000000000000011",--27698
"001001111100000111111111111111111000",--27699
"000111000000000000000111010110110001",--27700
"101000000011111000000001000000000000",--27701
"101001000000000000010000000000000101",--27702
"000111000000000000000111010110101010",--27703
"001101111100000111111111111111111000",--27704
"101110000001111000000001100000000000",--27705
"001001111100000000011111111111111000",--27706
"101001000000000000010000000000000011",--27707
"001001111100000111111111111111110111",--27708
"000111000000000000000111010110110001",--27709
"001101111100000000101111111111111000",--27710
"001001000100000000010000000000000001",--27711
"101001000000000000010000000000000011",--27712
"101110000001111000000001100000000000",--27713
"000111000000000000000111010110110001",--27714
"001101111100000000101111111111111000",--27715
"001001000100000000010000000000000010",--27716
"101001000000000000010000000000000011",--27717
"101110000001111000000001100000000000",--27718
"000111000000000000000111010110110001",--27719
"001101111100000000101111111111111000",--27720
"001001000100000000010000000000000011",--27721
"101001000000000000010000000000000011",--27722
"101110000001111000000001100000000000",--27723
"000111000000000000000111010110110001",--27724
"001101111100000000101111111111111000",--27725
"001001000100000000010000000000000100",--27726
"101000111011111000000000100000000000",--27727
"101001111010000111010000000000001000",--27728
"001001000010000000100000000000000111",--27729
"001101111100000000101111111111111001",--27730
"001001000010000000100000000000000110",--27731
"001101111100000000101111111111111010",--27732
"001001000010000000100000000000000101",--27733
"001101111100000000101111111111111011",--27734
"001001000010000000100000000000000100",--27735
"001101111100000000101111111111111100",--27736
"001001000010000000100000000000000011",--27737
"001101111100000000101111111111111101",--27738
"001001000010000000100000000000000010",--27739
"001101111100000000101111111111111110",--27740
"001001000010000000100000000000000001",--27741
"001101111100000000101111111111111111",--27742
"001001000010000000100000000000000000",--27743
"101000000011111000000001000000000000",--27744
"001101111100000000010000000000000000",--27745
"000111000000000000000111010110101010",--27746
"001101111100000111111111111111110111",--27747
"001101000000000000100000000100011011",--27748
"101001000100010000100000000000000010",--27749
"010111000100000000001111100000000000",--27750
"000101000000000000000110101100011000",--27751
"011011000011000001010000001000101000",--27752
"111110001000001001000001100000000000",--27753
"101111001001110001000011110111001100",--27754
"101111001001100001001100110011001101",--27755
"111110000110000001000001100000000000",--27756
"111110000110100000000001100000000000",--27757
"111110000110011000000010000000000000",--27758
"010110001001000000010000000000000010",--27759
"101001000000000001000000000000000001",--27760
"000101000000000000000110110001110111",--27761
"011010001001000000100000000000000010",--27762
"101001000000000001001111111111111111",--27763
"000101000000000000000110110001110111",--27764
"101000000001111000000010000000000000",--27765
"000101000000000000000110110001111000",--27766
"111110001000011000000010000000000000",--27767
"111110001000001001000011100000000000",--27768
"101111000001110010000100001011110010",--27769
"111110010000001001110100000000000000",--27770
"101111010011110010010011110100110010",--27771
"101111010011100010010001011001000011",--27772
"111110010000001010010100000000000000",--27773
"101111000001110010010100001011001000",--27774
"111110010010001001110100100000000000",--27775
"101111000001110010100100000110101000",--27776
"111110010100000010000100000000000000",--27777
"111110010000011000000100000000000000",--27778
"111110010010001010000100000000000000",--27779
"101111000001110010010100001010100010",--27780
"111110010010001001110100100000000000",--27781
"101111000001110010100100000110011000",--27782
"111110010100000010000100000000000000",--27783
"111110010000011000000100000000000000",--27784
"111110010010001010000100000000000000",--27785
"101111000001110010010100001010000000",--27786
"111110010010001001110100100000000000",--27787
"101111000001110010100100000110001000",--27788
"111110010100000010000100000000000000",--27789
"111110010000011000000100000000000000",--27790
"111110010010001010000100000000000000",--27791
"101111000001110010010100001001000100",--27792
"111110010010001001110100100000000000",--27793
"101111000001110010100100000101110000",--27794
"111110010100000010000100000000000000",--27795
"111110010000011000000100000000000000",--27796
"111110010010001010000100000000000000",--27797
"101111000001110010010100001000010000",--27798
"111110010010001001110100100000000000",--27799
"101111000001110010100100000101010000",--27800
"111110010100000010000100000000000000",--27801
"111110010000011000000100000000000000",--27802
"111110010010001010000100000000000000",--27803
"101111000001110010010100000111001000",--27804
"111110010010001001110100100000000000",--27805
"101111000001110010100100000100110000",--27806
"111110010100000010000100000000000000",--27807
"111110010000011000000100000000000000",--27808
"111110010010001010000100000000000000",--27809
"101111000001110010010100000110000000",--27810
"111110010010001001110100100000000000",--27811
"101111000001110010100100000100010000",--27812
"111110010100000010000100000000000000",--27813
"111110010000011000000100000000000000",--27814
"111110010010001010000100000000000000",--27815
"101111000001110010010100000100010000",--27816
"111110010010001001110100100000000000",--27817
"101111000001110010100100000011100000",--27818
"111110010100000010000100000000000000",--27819
"111110010000011000000100000000000000",--27820
"111110010010001010000100000000000000",--27821
"101111000001110010010100000010000000",--27822
"111110010010001001110100100000000000",--27823
"101111000001110010100100000010100000",--27824
"111110010100000010000100000000000000",--27825
"111110010000011000000100000000000000",--27826
"111110010010001010000100000000000000",--27827
"101111000001110010010100000001000000",--27828
"111110010010000010000100000000000000",--27829
"111110010000011000000100000000000000",--27830
"111110001110001010000011100000000000",--27831
"111110001110000000010011100000000000",--27832
"111110001110011000000011100000000000",--27833
"111110001000001001110010000000000000",--27834
"010100001001000000000000000000000100",--27835
"101111001111110001110011111111001001",--27836
"101111001111100001110000111111011010",--27837
"111110001110010001000010000000000000",--27838
"000101000000000000000110110011000100",--27839
"011000001001000000000000000000000011",--27840
"101111001111110001111011111111001001",--27841
"101111001111100001110000111111011010",--27842
"111110001110010001000010000000000000",--27843
"111110001000001001010010000000000000",--27844
"111110001000001001000011100000000000",--27845
"101111000001110010000100000011100000",--27846
"101111010011110010010011110111100011",--27847
"101111010011100010011000111000111001",--27848
"111110001110001010010100100000000000",--27849
"101111000001110010100100000010100000",--27850
"111110010000010010010100000000000000",--27851
"111110010000011000000100000000000000",--27852
"111110001110001010000100000000000000",--27853
"101111000001110010010100000001000000",--27854
"111110010100010010000100000000000000",--27855
"111110010000011000000100000000000000",--27856
"111110001110001010000100000000000000",--27857
"111110010010010010000100000000000000",--27858
"111110010000011000000100000000000000",--27859
"111110001110001010000011100000000000",--27860
"111110001110010000010011100000000010",--27861
"111110001110011000000011100000000000",--27862
"111110001000001001110010000000000000",--27863
"111110001000001000110001100000000000",--27864
"101001000010000000010000000000000001",--27865
"111110000110001000110010000000000000",--27866
"101111001111110001110011110111001100",--27867
"101111001111100001111100110011001101",--27868
"111110001000000001110010000000000000",--27869
"111110001000100000000010000000000000",--27870
"111110001000011000000011100000000000",--27871
"010110001111000000010000000000000010",--27872
"101001000000000001000000000000000001",--27873
"000101000000000000000110110011101000",--27874
"011010001111000000100000000000000010",--27875
"101001000000000001001111111111111111",--27876
"000101000000000000000110110011101000",--27877
"101000000001111000000010000000000000",--27878
"000101000000000000000110110011101001",--27879
"111110001110011000000011100000000000",--27880
"111110001110001001110100000000000000",--27881
"101111000001110010010100001011110010",--27882
"111110010010001010000100100000000000",--27883
"101111010101110010100011110100110010",--27884
"101111010101100010100001011001000011",--27885
"111110010010001010100100100000000000",--27886
"101111000001110010100100001011001000",--27887
"111110010100001010000101000000000000",--27888
"101111000001110010110100000110101000",--27889
"111110010110000010010100100000000000",--27890
"111110010010011000000100100000000000",--27891
"111110010100001010010100100000000000",--27892
"101111000001110010100100001010100010",--27893
"111110010100001010000101000000000000",--27894
"101111000001110010110100000110011000",--27895
"111110010110000010010100100000000000",--27896
"111110010010011000000100100000000000",--27897
"111110010100001010010100100000000000",--27898
"101111000001110010100100001010000000",--27899
"111110010100001010000101000000000000",--27900
"101111000001110010110100000110001000",--27901
"111110010110000010010100100000000000",--27902
"111110010010011000000100100000000000",--27903
"111110010100001010010100100000000000",--27904
"101111000001110010100100001001000100",--27905
"111110010100001010000101000000000000",--27906
"101111000001110010110100000101110000",--27907
"111110010110000010010100100000000000",--27908
"111110010010011000000100100000000000",--27909
"111110010100001010010100100000000000",--27910
"101111000001110010100100001000010000",--27911
"111110010100001010000101000000000000",--27912
"101111000001110010110100000101010000",--27913
"111110010110000010010100100000000000",--27914
"111110010010011000000100100000000000",--27915
"111110010100001010010100100000000000",--27916
"101111000001110010100100000111001000",--27917
"111110010100001010000101000000000000",--27918
"101111000001110010110100000100110000",--27919
"111110010110000010010100100000000000",--27920
"111110010010011000000100100000000000",--27921
"111110010100001010010100100000000000",--27922
"101111000001110010100100000110000000",--27923
"111110010100001010000101000000000000",--27924
"101111000001110010110100000100010000",--27925
"111110010110000010010100100000000000",--27926
"111110010010011000000100100000000000",--27927
"111110010100001010010100100000000000",--27928
"101111000001110010100100000100010000",--27929
"111110010100001010000101000000000000",--27930
"101111000001110010110100000011100000",--27931
"111110010110000010010100100000000000",--27932
"111110010010011000000100100000000000",--27933
"111110010100001010010100100000000000",--27934
"101111000001110010100100000010000000",--27935
"111110010100001010000101000000000000",--27936
"101111000001110010110100000010100000",--27937
"111110010110000010010100100000000000",--27938
"111110010010011000000100100000000000",--27939
"111110010100001010010100100000000000",--27940
"101111000001110010100100000001000000",--27941
"111110010100000010010100100000000000",--27942
"111110010010011000000100100000000000",--27943
"111110010000001010010100000000000000",--27944
"111110010000000000010100000000000000",--27945
"111110010000011000000100000000000000",--27946
"111110001110001010000011100000000000",--27947
"010100001001000000000000000000000100",--27948
"101111010001110010000011111111001001",--27949
"101111010001100010000000111111011010",--27950
"111110010000010001110011100000000000",--27951
"000101000000000000000110110100110101",--27952
"011000001001000000000000000000000011",--27953
"101111010001110010001011111111001001",--27954
"101111010001100010000000111111011010",--27955
"111110010000010001110011100000000000",--27956
"111110001110001001100011100000000000",--27957
"111110001110001001110100000000000000",--27958
"101111000001110010010100000011100000",--27959
"101111010101110010100011110111100011",--27960
"101111010101100010101000111000111001",--27961
"111110010000001010100101000000000000",--27962
"101111000001110010110100000010100000",--27963
"111110010010010010100100100000000000",--27964
"111110010010011000000100100000000000",--27965
"111110010000001010010100100000000000",--27966
"101111000001110010100100000001000000",--27967
"111110010110010010010100100000000000",--27968
"111110010010011000000100100000000000",--27969
"111110010000001010010100100000000000",--27970
"111110010100010010010100100000000000",--27971
"111110010010011000000100100000000000",--27972
"111110010000001010010100000000000000",--27973
"111110010000010000010100000000000010",--27974
"111110010000011000000100000000000000",--27975
"111110001110001010000011100000000000",--27976
"111110001110001001000010000000000000",--27977
"011011000011000001010000000100001110",--27978
"111110001000001001000001100000000000",--27979
"101111001001110001000011110111001100",--27980
"101111001001100001001100110011001101",--27981
"111110000110000001000001100000000000",--27982
"111110000110100000000001100000000000",--27983
"111110000110011000000010000000000000",--27984
"010110001001000000010000000000000010",--27985
"101001000000000001000000000000000001",--27986
"000101000000000000000110110101011001",--27987
"011010001001000000100000000000000010",--27988
"101001000000000001001111111111111111",--27989
"000101000000000000000110110101011001",--27990
"101000000001111000000010000000000000",--27991
"000101000000000000000110110101011010",--27992
"111110001000011000000010000000000000",--27993
"111110001000001001000011100000000000",--27994
"101111000001110010000100001011110010",--27995
"111110010000001001110100000000000000",--27996
"101111010011110010010011110100110010",--27997
"101111010011100010010001011001000011",--27998
"111110010000001010010100000000000000",--27999
"101111000001110010010100001011001000",--28000
"111110010010001001110100100000000000",--28001
"101111000001110010100100000110101000",--28002
"111110010100000010000100000000000000",--28003
"111110010000011000000100000000000000",--28004
"111110010010001010000100000000000000",--28005
"101111000001110010010100001010100010",--28006
"111110010010001001110100100000000000",--28007
"101111000001110010100100000110011000",--28008
"111110010100000010000100000000000000",--28009
"111110010000011000000100000000000000",--28010
"111110010010001010000100000000000000",--28011
"101111000001110010010100001010000000",--28012
"111110010010001001110100100000000000",--28013
"101111000001110010100100000110001000",--28014
"111110010100000010000100000000000000",--28015
"111110010000011000000100000000000000",--28016
"111110010010001010000100000000000000",--28017
"101111000001110010010100001001000100",--28018
"111110010010001001110100100000000000",--28019
"101111000001110010100100000101110000",--28020
"111110010100000010000100000000000000",--28021
"111110010000011000000100000000000000",--28022
"111110010010001010000100000000000000",--28023
"101111000001110010010100001000010000",--28024
"111110010010001001110100100000000000",--28025
"101111000001110010100100000101010000",--28026
"111110010100000010000100000000000000",--28027
"111110010000011000000100000000000000",--28028
"111110010010001010000100000000000000",--28029
"101111000001110010010100000111001000",--28030
"111110010010001001110100100000000000",--28031
"101111000001110010100100000100110000",--28032
"111110010100000010000100000000000000",--28033
"111110010000011000000100000000000000",--28034
"111110010010001010000100000000000000",--28035
"101111000001110010010100000110000000",--28036
"111110010010001001110100100000000000",--28037
"101111000001110010100100000100010000",--28038
"111110010100000010000100000000000000",--28039
"111110010000011000000100000000000000",--28040
"111110010010001010000100000000000000",--28041
"101111000001110010010100000100010000",--28042
"111110010010001001110100100000000000",--28043
"101111000001110010100100000011100000",--28044
"111110010100000010000100000000000000",--28045
"111110010000011000000100000000000000",--28046
"111110010010001010000100000000000000",--28047
"101111000001110010010100000010000000",--28048
"111110010010001001110100100000000000",--28049
"101111000001110010100100000010100000",--28050
"111110010100000010000100000000000000",--28051
"111110010000011000000100000000000000",--28052
"111110010010001010000100000000000000",--28053
"101111000001110010100100000001000000",--28054
"111110010100000010000100000000000000",--28055
"111110010000011000000100000000000000",--28056
"111110001110001010000100000000000000",--28057
"001001111100000000110000000000000000",--28058
"001001111100000000101111111111111111",--28059
"001011111100000001101111111111111110",--28060
"001001111100000000011111111111111101",--28061
"001011111100000000111111111111111100",--28062
"001011111100000001011111111111111011",--28063
"001001111100000001001111111111111010",--28064
"001011111100000001001111111111111001",--28065
"101110010001111000000010100000000000",--28066
"101110001111111000000010000000000000",--28067
"101110000001111000000001100000000000",--28068
"001001111100000111111111111111111000",--28069
"101001111100010111100000000000001001",--28070
"000111000000000000000000001101001100",--28071
"101001111100000111100000000000001001",--28072
"001101111100000111111111111111111000",--28073
"111110000110000000010001100000000000",--28074
"111110000110011000000001100000000000",--28075
"001111111100000001001111111111111001",--28076
"111110001000001000110001100000000000",--28077
"001101111100000000011111111111111010",--28078
"010100000011000000000000000000000100",--28079
"101111001001110001000011111111001001",--28080
"101111001001100001000000111111011010",--28081
"111110001000010000110001100000000000",--28082
"000101000000000000000110110110111000",--28083
"011000000011000000000000000000000011",--28084
"101111001001110001001011111111001001",--28085
"101111001001100001000000111111011010",--28086
"111110001000010000110001100000000000",--28087
"001111111100000001001111111111111011",--28088
"111110000110001001000001100000000000",--28089
"111110000110001000110010100000000000",--28090
"101111000001110001100100000011100000",--28091
"101111001111110001110011110111100011",--28092
"101111001111100001111000111000111001",--28093
"111110001010001001110011100000000000",--28094
"101111000001110010000100000010100000",--28095
"111110001100010001110011000000000000",--28096
"111110001100011000000011000000000000",--28097
"111110001010001001100011000000000000",--28098
"101111000001110001110100000001000000",--28099
"111110010000010001100011000000000000",--28100
"111110001100011000000011000000000000",--28101
"111110001010001001100011000000000000",--28102
"111110001110010001100011000000000000",--28103
"111110001100011000000011000000000000",--28104
"111110001010001001100010100000000000",--28105
"111110001010010000010010100000000010",--28106
"111110001010011000000010100000000000",--28107
"111110000110001001010001100000000000",--28108
"001111111100000001011111111111111100",--28109
"111110000110001001010001100000000000",--28110
"001101111100000000011111111111111101",--28111
"101001000010000000010000000000000001",--28112
"111110000110001000110010100000000000",--28113
"101111001101110001100011110111001100",--28114
"101111001101100001101100110011001101",--28115
"111110001010000001100010100000000000",--28116
"111110001010100000000010100000000000",--28117
"111110001010011000000011000000000000",--28118
"010110001101000000010000000000000010",--28119
"101001000000000000100000000000000001",--28120
"000101000000000000000110110111011111",--28121
"011010001101000000100000000000000010",--28122
"101001000000000000101111111111111111",--28123
"000101000000000000000110110111011111",--28124
"101000000001111000000001000000000000",--28125
"000101000000000000000110110111100000",--28126
"111110001100011000000011000000000000",--28127
"111110001100001001100011100000000000",--28128
"101111000001110010000100001011110010",--28129
"111110010000001001110100000000000000",--28130
"101111010011110010010011110100110010",--28131
"101111010011100010010001011001000011",--28132
"111110010000001010010100000000000000",--28133
"101111000001110010010100001011001000",--28134
"111110010010001001110100100000000000",--28135
"101111000001110010100100000110101000",--28136
"111110010100000010000100000000000000",--28137
"111110010000011000000100000000000000",--28138
"111110010010001010000100000000000000",--28139
"101111000001110010010100001010100010",--28140
"111110010010001001110100100000000000",--28141
"101111000001110010100100000110011000",--28142
"111110010100000010000100000000000000",--28143
"111110010000011000000100000000000000",--28144
"111110010010001010000100000000000000",--28145
"101111000001110010010100001010000000",--28146
"111110010010001001110100100000000000",--28147
"101111000001110010100100000110001000",--28148
"111110010100000010000100000000000000",--28149
"111110010000011000000100000000000000",--28150
"111110010010001010000100000000000000",--28151
"101111000001110010010100001001000100",--28152
"111110010010001001110100100000000000",--28153
"101111000001110010100100000101110000",--28154
"111110010100000010000100000000000000",--28155
"111110010000011000000100000000000000",--28156
"111110010010001010000100000000000000",--28157
"101111000001110010010100001000010000",--28158
"111110010010001001110100100000000000",--28159
"101111000001110010100100000101010000",--28160
"111110010100000010000100000000000000",--28161
"111110010000011000000100000000000000",--28162
"111110010010001010000100000000000000",--28163
"101111000001110010010100000111001000",--28164
"111110010010001001110100100000000000",--28165
"101111000001110010100100000100110000",--28166
"111110010100000010000100000000000000",--28167
"111110010000011000000100000000000000",--28168
"111110010010001010000100000000000000",--28169
"101111000001110010010100000110000000",--28170
"111110010010001001110100100000000000",--28171
"101111000001110010100100000100010000",--28172
"111110010100000010000100000000000000",--28173
"111110010000011000000100000000000000",--28174
"111110010010001010000100000000000000",--28175
"101111000001110010010100000100010000",--28176
"111110010010001001110100100000000000",--28177
"101111000001110010100100000011100000",--28178
"111110010100000010000100000000000000",--28179
"111110010000011000000100000000000000",--28180
"111110010010001010000100000000000000",--28181
"101111000001110010010100000010000000",--28182
"111110010010001001110100100000000000",--28183
"101111000001110010100100000010100000",--28184
"111110010100000010000100000000000000",--28185
"111110010000011000000100000000000000",--28186
"111110010010001010000100000000000000",--28187
"101111000001110010100100000001000000",--28188
"111110010100000010000100000000000000",--28189
"111110010000011000000100000000000000",--28190
"111110001110001010000100000000000000",--28191
"001011111100000000111111111111111000",--28192
"001001111100000000011111111111110111",--28193
"001011111100000001011111111111110110",--28194
"001001111100000000101111111111110101",--28195
"001011111100000001101111111111110100",--28196
"101110010001111000000010100000000000",--28197
"101110001111111000000010000000000000",--28198
"101110000001111000000001100000000000",--28199
"001001111100000111111111111111110011",--28200
"101001111100010111100000000000001110",--28201
"000111000000000000000000001101001100",--28202
"101001111100000111100000000000001110",--28203
"001101111100000111111111111111110011",--28204
"111110000110000000010001100000000000",--28205
"111110000110011000000001100000000000",--28206
"001111111100000001001111111111110100",--28207
"111110001000001000110001100000000000",--28208
"001101111100000000011111111111110101",--28209
"010100000011000000000000000000000100",--28210
"101111001001110001000011111111001001",--28211
"101111001001100001000000111111011010",--28212
"111110001000010000110001100000000000",--28213
"000101000000000000000110111000111011",--28214
"011000000011000000000000000000000011",--28215
"101111001001110001001011111111001001",--28216
"101111001001100001000000111111011010",--28217
"111110001000010000110001100000000000",--28218
"001111111100000001101111111111111110",--28219
"111110000110001001100001100000000000",--28220
"111110000110001000110010000000000000",--28221
"101111000001110001010100000011100000",--28222
"101111001111110001110011110111100011",--28223
"101111001111100001111000111000111001",--28224
"111110001000001001110011100000000000",--28225
"101111000001110010000100000010100000",--28226
"111110001010010001110010100000000000",--28227
"111110001010011000000010100000000000",--28228
"111110001000001001010010100000000000",--28229
"101111000001110001110100000001000000",--28230
"111110010000010001010010100000000000",--28231
"111110001010011000000010100000000000",--28232
"111110001000001001010010100000000000",--28233
"111110001110010001010010100000000000",--28234
"111110001010011000000010100000000000",--28235
"111110001000001001010010000000000000",--28236
"111110001000010000010010000000000010",--28237
"111110001000011000000010000000000000",--28238
"111110000110001001000001100000000000",--28239
"001111111100000001001111111111110110",--28240
"111110000110001001000010000000000000",--28241
"001111111100000000111111111111111000",--28242
"001111111100000001011111111111111011",--28243
"001101111100000000011111111111110111",--28244
"001101111100000000101111111111111111",--28245
"001101111100000000110000000000000000",--28246
"011011000011000001010000000000111001",--28247
"000101000000000000000110110001101001",--28248
"111110000110001000110010100000000000",--28249
"111110001000001001000011000000000000",--28250
"111110001010000001100010100000000000",--28251
"111110001010000000010010100000000000",--28252
"111110001010100000000010100000000000",--28253
"111110001010011000000011000000000000",--28254
"111110000110001001100001100000000000",--28255
"111110001010011000000011000000000000",--28256
"111110001000001001100010000000000000",--28257
"111110001010011000000010100000000000",--28258
"001101000100000000010000000011111110",--28259
"001100000010000000110001000000000000",--28260
"001101000100000000100000000000000000",--28261
"001011000100000000110000000000000000",--28262
"001011000100000001000000000000000001",--28263
"001011000100000001010000000000000010",--28264
"101001000110000000100000000000101000",--28265
"001100000010000000100001000000000000",--28266
"001101000100000000100000000000000000",--28267
"101110001001111000000011000000000010",--28268
"001011000100000000110000000000000000",--28269
"001011000100000001010000000000000001",--28270
"001011000100000001100000000000000010",--28271
"101001000110000000100000000001010000",--28272
"001100000010000000100001000000000000",--28273
"001101000100000000100000000000000000",--28274
"101110000111111000000011000000000010",--28275
"101110001001111000000011100000000010",--28276
"001011000100000001010000000000000000",--28277
"001011000100000001100000000000000001",--28278
"001011000100000001110000000000000010",--28279
"101001000110000000100000000000000001",--28280
"001100000010000000100001000000000000",--28281
"001101000100000000100000000000000000",--28282
"101110000111111000000011000000000010",--28283
"101110001001111000000011100000000010",--28284
"101110001011111000000100000000000010",--28285
"001011000100000001100000000000000000",--28286
"001011000100000001110000000000000001",--28287
"001011000100000010000000000000000010",--28288
"101001000110000000100000000000101001",--28289
"001100000010000000100001000000000000",--28290
"001101000100000000100000000000000000",--28291
"101110000111111000000011000000000010",--28292
"101110001011111000000011100000000010",--28293
"001011000100000001100000000000000000",--28294
"001011000100000001110000000000000001",--28295
"001011000100000001000000000000000010",--28296
"101001000110000000100000000001010001",--28297
"001100000010000000100000100000000000",--28298
"001101000010000000010000000000000000",--28299
"101110001011111000000010100000000010",--28300
"001011000010000001010000000000000000",--28301
"001011000010000000110000000000000001",--28302
"001011000010000001000000000000000010",--28303
"000100000000000000001111100000000000",--28304
"111110000110001000110010100000000000",--28305
"111110001000001001000011000000000000",--28306
"111110001010000001100010100000000000",--28307
"111110001010000000010010100000000000",--28308
"111110001010100000000010100000000000",--28309
"111110001010011000000011000000000000",--28310
"111110000110001001100001100000000000",--28311
"111110001010011000000011000000000000",--28312
"111110001000001001100010000000000000",--28313
"111110001010011000000010100000000000",--28314
"001101000100000000010000000011111110",--28315
"001100000010000000110001000000000000",--28316
"001101000100000000100000000000000000",--28317
"001011000100000000110000000000000000",--28318
"001011000100000001000000000000000001",--28319
"001011000100000001010000000000000010",--28320
"101001000110000000100000000000101000",--28321
"001100000010000000100001000000000000",--28322
"001101000100000000100000000000000000",--28323
"101110001001111000000011000000000010",--28324
"001011000100000000110000000000000000",--28325
"001011000100000001010000000000000001",--28326
"001011000100000001100000000000000010",--28327
"101001000110000000100000000001010000",--28328
"001100000010000000100001000000000000",--28329
"001101000100000000100000000000000000",--28330
"101110000111111000000011000000000010",--28331
"101110001001111000000011100000000010",--28332
"001011000100000001010000000000000000",--28333
"001011000100000001100000000000000001",--28334
"001011000100000001110000000000000010",--28335
"101001000110000000100000000000000001",--28336
"001100000010000000100001000000000000",--28337
"001101000100000000100000000000000000",--28338
"101110000111111000000011000000000010",--28339
"101110001001111000000011100000000010",--28340
"101110001011111000000100000000000010",--28341
"001011000100000001100000000000000000",--28342
"001011000100000001110000000000000001",--28343
"001011000100000010000000000000000010",--28344
"101001000110000000100000000000101001",--28345
"001100000010000000100001000000000000",--28346
"001101000100000000100000000000000000",--28347
"101110000111111000000011000000000010",--28348
"101110001011111000000011100000000010",--28349
"001011000100000001100000000000000000",--28350
"001011000100000001110000000000000001",--28351
"001011000100000001000000000000000010",--28352
"101001000110000000100000000001010001",--28353
"001100000010000000100000100000000000",--28354
"001101000010000000010000000000000000",--28355
"101110001011111000000010100000000010",--28356
"001011000010000001010000000000000000",--28357
"001011000010000000110000000000000001",--28358
"001011000010000001000000000000000010",--28359
"000100000000000000001111100000000000",--28360
"010111000010000000001111100000000000",--28361
"101010000011101000000010000000000000",--28362
"101111001011110001010011111001001100",--28363
"101111001011100001011100110011001101",--28364
"111110001000001001010010000000000000",--28365
"101111001011110001010011111101100110",--28366
"101111001011100001010110011001100110",--28367
"111110001000010001010010000000000000",--28368
"101111001011110001010011111010100001",--28369
"101111001011100001011110100010011001",--28370
"101111001101110001100011111010100001",--28371
"101111001101100001101110100010011000",--28372
"101111001111110001110011110111001100",--28373
"101111001111100001111100110011000101",--28374
"101111010011110010010011110100000101",--28375
"101111010011100010010001001001010001",--28376
"001001111100000000010000000000000000",--28377
"001001111100000000111111111111111111",--28378
"001001111100000000101111111111111110",--28379
"001011111100000000111111111111111101",--28380
"001011111100000001011111111111111100",--28381
"001011111100000001001111111111111011",--28382
"001011111100000001101111111111111010",--28383
"101110010011111000000010100000000000",--28384
"101110001111111000000010000000000000",--28385
"101110000001111000000001100000000000",--28386
"001001111100000111111111111111111001",--28387
"101001111100010111100000000000001000",--28388
"000111000000000000000000001101001100",--28389
"101001111100000111100000000000001000",--28390
"001101111100000111111111111111111001",--28391
"111110000110000000010001100000000000",--28392
"111110000110011000000001100000000000",--28393
"001111111100000001001111111111111010",--28394
"111110001000001000110001100000000000",--28395
"101111001001110001000011111111001001",--28396
"101111001001100001000000111111011010",--28397
"111110001000010000110001100000000000",--28398
"001111111100000001001111111111111011",--28399
"111110000110001001000001100000000000",--28400
"111110000110001000110010100000000000",--28401
"101111000001110001100100000011100000",--28402
"101111001111110001110011110111100011",--28403
"101111001111100001111000111000111001",--28404
"111110001010001001110011100000000000",--28405
"101111000001110010000100000010100000",--28406
"111110001100010001110011000000000000",--28407
"111110001100011000000011000000000000",--28408
"111110001010001001100011000000000000",--28409
"101111000001110001110100000001000000",--28410
"111110010000010001100011000000000000",--28411
"111110001100011000000011000000000000",--28412
"111110001010001001100011000000000000",--28413
"111110001110010001100011000000000000",--28414
"111110001100011000000011000000000000",--28415
"111110001010001001100010100000000000",--28416
"111110001010010000010010100000000010",--28417
"111110001010011000000010100000000000",--28418
"111110000110001001010001100000000000",--28419
"001111111100000001011111111111111100",--28420
"111110000110001001010001100000000000",--28421
"101001000000000000010000000000000001",--28422
"111110000110001000110010100000000000",--28423
"101111001101110001100011110111001100",--28424
"101111001101100001101100110011001101",--28425
"111110001010000001100010100000000000",--28426
"111110001010100000000010100000000000",--28427
"111110001010011000000011000000000000",--28428
"010110001101000000010000000000000010",--28429
"101001000000000000100000000000000001",--28430
"000101000000000000000110111100010101",--28431
"011010001101000000100000000000000010",--28432
"101001000000000000101111111111111111",--28433
"000101000000000000000110111100010101",--28434
"101000000001111000000001000000000000",--28435
"000101000000000000000110111100010110",--28436
"111110001100011000000011000000000000",--28437
"111110001100001001100011100000000000",--28438
"101111000001110010000100001011110010",--28439
"111110010000001001110100000000000000",--28440
"101111010011110010010011110100110010",--28441
"101111010011100010010001011001000011",--28442
"111110010000001010010100000000000000",--28443
"101111000001110010010100001011001000",--28444
"111110010010001001110100100000000000",--28445
"101111000001110010100100000110101000",--28446
"111110010100000010000100000000000000",--28447
"111110010000011000000100000000000000",--28448
"111110010010001010000100000000000000",--28449
"101111000001110010010100001010100010",--28450
"111110010010001001110100100000000000",--28451
"101111000001110010100100000110011000",--28452
"111110010100000010000100000000000000",--28453
"111110010000011000000100000000000000",--28454
"111110010010001010000100000000000000",--28455
"101111000001110010010100001010000000",--28456
"111110010010001001110100100000000000",--28457
"101111000001110010100100000110001000",--28458
"111110010100000010000100000000000000",--28459
"111110010000011000000100000000000000",--28460
"111110010010001010000100000000000000",--28461
"101111000001110010010100001001000100",--28462
"111110010010001001110100100000000000",--28463
"101111000001110010100100000101110000",--28464
"111110010100000010000100000000000000",--28465
"111110010000011000000100000000000000",--28466
"111110010010001010000100000000000000",--28467
"101111000001110010010100001000010000",--28468
"111110010010001001110100100000000000",--28469
"101111000001110010100100000101010000",--28470
"111110010100000010000100000000000000",--28471
"111110010000011000000100000000000000",--28472
"111110010010001010000100000000000000",--28473
"101111000001110010010100000111001000",--28474
"111110010010001001110100100000000000",--28475
"101111000001110010100100000100110000",--28476
"111110010100000010000100000000000000",--28477
"111110010000011000000100000000000000",--28478
"111110010010001010000100000000000000",--28479
"101111000001110010010100000110000000",--28480
"111110010010001001110100100000000000",--28481
"101111000001110010100100000100010000",--28482
"111110010100000010000100000000000000",--28483
"111110010000011000000100000000000000",--28484
"111110010010001010000100000000000000",--28485
"101111000001110010010100000100010000",--28486
"111110010010001001110100100000000000",--28487
"101111000001110010100100000011100000",--28488
"111110010100000010000100000000000000",--28489
"111110010000011000000100000000000000",--28490
"111110010010001010000100000000000000",--28491
"101111000001110010010100000010000000",--28492
"111110010010001001110100100000000000",--28493
"101111000001110010100100000010100000",--28494
"111110010100000010000100000000000000",--28495
"111110010000011000000100000000000000",--28496
"111110010010001010000100000000000000",--28497
"101111000001110010100100000001000000",--28498
"111110010100000010000100000000000000",--28499
"111110010000011000000100000000000000",--28500
"111110001110001010000100000000000000",--28501
"001011111100000000111111111111111001",--28502
"001001111100000000011111111111111000",--28503
"001011111100000001011111111111110111",--28504
"001001111100000000101111111111110110",--28505
"001011111100000001101111111111110101",--28506
"101110010001111000000010100000000000",--28507
"101110001111111000000010000000000000",--28508
"101110000001111000000001100000000000",--28509
"001001111100000111111111111111110100",--28510
"101001111100010111100000000000001101",--28511
"000111000000000000000000001101001100",--28512
"101001111100000111100000000000001101",--28513
"001101111100000111111111111111110100",--28514
"111110000110000000010001100000000000",--28515
"111110000110011000000001100000000000",--28516
"001111111100000001001111111111110101",--28517
"111110001000001000110001100000000000",--28518
"001101111100000000011111111111110110",--28519
"010100000011000000000000000000000100",--28520
"101111001001110001000011111111001001",--28521
"101111001001100001000000111111011010",--28522
"111110001000010000110001100000000000",--28523
"000101000000000000000110111101110001",--28524
"011000000011000000000000000000000011",--28525
"101111001001110001001011111111001001",--28526
"101111001001100001000000111111011010",--28527
"111110001000010000110001100000000000",--28528
"001111111100000001101111111111111101",--28529
"111110000110001001100001100000000000",--28530
"111110000110001000110010000000000000",--28531
"101111000001110001010100000011100000",--28532
"101111001111110001110011110111100011",--28533
"101111001111100001111000111000111001",--28534
"111110001000001001110011100000000000",--28535
"101111000001110010000100000010100000",--28536
"111110001010010001110010100000000000",--28537
"111110001010011000000010100000000000",--28538
"111110001000001001010010100000000000",--28539
"101111000001110001110100000001000000",--28540
"111110010000010001010010100000000000",--28541
"111110001010011000000010100000000000",--28542
"111110001000001001010010100000000000",--28543
"111110001110010001010010100000000000",--28544
"111110001010011000000010100000000000",--28545
"111110001000001001010010000000000000",--28546
"111110001000010000010010000000000010",--28547
"111110001000011000000010000000000000",--28548
"111110000110001001000001100000000000",--28549
"001111111100000001001111111111110111",--28550
"111110000110001001000010000000000000",--28551
"001111111100000000111111111111111001",--28552
"001111111100000001011111111111111011",--28553
"001101111100000000011111111111111000",--28554
"001101111100000000101111111111111110",--28555
"001101111100000000111111111111111111",--28556
"001001111100000111111111111111110100",--28557
"101001111100010111100000000000001101",--28558
"000111000000000000000110110001101000",--28559
"101001111100000111100000000000001101",--28560
"001101111100000111111111111111110100",--28561
"001101111100000000011111111111111111",--28562
"101001000010000000100000000000000010",--28563
"001101111100000000110000000000000000",--28564
"101010000111101000000001100000000000",--28565
"101111001001110001000011111001001100",--28566
"101111001001100001001100110011001101",--28567
"111110000110001001000001100000000000",--28568
"101111001001110001000011110111001100",--28569
"101111001001100001001100110011001101",--28570
"111110000110000001000001100000000000",--28571
"101111001001110001000011111010100001",--28572
"101111001001100001001110100010011001",--28573
"101111001011110001010011111010100001",--28574
"101111001011100001011110100010011000",--28575
"101111001101110001100011110111001100",--28576
"101111001101100001101100110011000101",--28577
"101111010001110010000011110100000101",--28578
"101111010001100010000001001001010001",--28579
"001001111100000000101111111111110100",--28580
"001011111100000001001111111111110011",--28581
"001011111100000000111111111111110010",--28582
"001011111100000001011111111111110001",--28583
"101110010001111000000010100000000000",--28584
"101110001101111000000010000000000000",--28585
"101110000001111000000001100000000000",--28586
"001001111100000111111111111111110000",--28587
"101001111100010111100000000000010001",--28588
"000111000000000000000000001101001100",--28589
"101001111100000111100000000000010001",--28590
"001101111100000111111111111111110000",--28591
"111110000110000000010001100000000000",--28592
"111110000110011000000001100000000000",--28593
"001111111100000001001111111111110001",--28594
"111110001000001000110001100000000000",--28595
"101111001001110001000011111111001001",--28596
"101111001001100001000000111111011010",--28597
"111110001000010000110001100000000000",--28598
"001111111100000001001111111111110010",--28599
"111110000110001001000001100000000000",--28600
"111110000110001000110010100000000000",--28601
"101111000001110001100100000011100000",--28602
"101111001111110001110011110111100011",--28603
"101111001111100001111000111000111001",--28604
"111110001010001001110011100000000000",--28605
"101111000001110010000100000010100000",--28606
"111110001100010001110011000000000000",--28607
"111110001100011000000011000000000000",--28608
"111110001010001001100011000000000000",--28609
"101111000001110001110100000001000000",--28610
"111110010000010001100011000000000000",--28611
"111110001100011000000011000000000000",--28612
"111110001010001001100011000000000000",--28613
"111110001110010001100011000000000000",--28614
"111110001100011000000011000000000000",--28615
"111110001010001001100010100000000000",--28616
"111110001010010000010010100000000010",--28617
"111110001010011000000010100000000000",--28618
"111110000110001001010001100000000000",--28619
"001111111100000001011111111111110011",--28620
"111110000110001001010001100000000000",--28621
"101001000000000000010000000000000001",--28622
"111110000110001000110010100000000000",--28623
"101111001101110001100011110111001100",--28624
"101111001101100001101100110011001101",--28625
"111110001010000001100010100000000000",--28626
"111110001010100000000010100000000000",--28627
"111110001010011000000011000000000000",--28628
"010110001101000000010000000000000010",--28629
"101001000000000000100000000000000001",--28630
"000101000000000000000110111111011101",--28631
"011010001101000000100000000000000010",--28632
"101001000000000000101111111111111111",--28633
"000101000000000000000110111111011101",--28634
"101000000001111000000001000000000000",--28635
"000101000000000000000110111111011110",--28636
"111110001100011000000011000000000000",--28637
"111110001100001001100011100000000000",--28638
"101111000001110010000100001011110010",--28639
"111110010000001001110100000000000000",--28640
"101111010011110010010011110100110010",--28641
"101111010011100010010001011001000011",--28642
"111110010000001010010100000000000000",--28643
"101111000001110010010100001011001000",--28644
"111110010010001001110100100000000000",--28645
"101111000001110010100100000110101000",--28646
"111110010100000010000100000000000000",--28647
"111110010000011000000100000000000000",--28648
"111110010010001010000100000000000000",--28649
"101111000001110010010100001010100010",--28650
"111110010010001001110100100000000000",--28651
"101111000001110010100100000110011000",--28652
"111110010100000010000100000000000000",--28653
"111110010000011000000100000000000000",--28654
"111110010010001010000100000000000000",--28655
"101111000001110010010100001010000000",--28656
"111110010010001001110100100000000000",--28657
"101111000001110010100100000110001000",--28658
"111110010100000010000100000000000000",--28659
"111110010000011000000100000000000000",--28660
"111110010010001010000100000000000000",--28661
"101111000001110010010100001001000100",--28662
"111110010010001001110100100000000000",--28663
"101111000001110010100100000101110000",--28664
"111110010100000010000100000000000000",--28665
"111110010000011000000100000000000000",--28666
"111110010010001010000100000000000000",--28667
"101111000001110010010100001000010000",--28668
"111110010010001001110100100000000000",--28669
"101111000001110010100100000101010000",--28670
"111110010100000010000100000000000000",--28671
"111110010000011000000100000000000000",--28672
"111110010010001010000100000000000000",--28673
"101111000001110010010100000111001000",--28674
"111110010010001001110100100000000000",--28675
"101111000001110010100100000100110000",--28676
"111110010100000010000100000000000000",--28677
"111110010000011000000100000000000000",--28678
"111110010010001010000100000000000000",--28679
"101111000001110010010100000110000000",--28680
"111110010010001001110100100000000000",--28681
"101111000001110010100100000100010000",--28682
"111110010100000010000100000000000000",--28683
"111110010000011000000100000000000000",--28684
"111110010010001010000100000000000000",--28685
"101111000001110010010100000100010000",--28686
"111110010010001001110100100000000000",--28687
"101111000001110010100100000011100000",--28688
"111110010100000010000100000000000000",--28689
"111110010000011000000100000000000000",--28690
"111110010010001010000100000000000000",--28691
"101111000001110010010100000010000000",--28692
"111110010010001001110100100000000000",--28693
"101111000001110010100100000010100000",--28694
"111110010100000010000100000000000000",--28695
"111110010000011000000100000000000000",--28696
"111110010010001010000100000000000000",--28697
"101111000001110010100100000001000000",--28698
"111110010100000010000100000000000000",--28699
"111110010000011000000100000000000000",--28700
"111110001110001010000100000000000000",--28701
"001011111100000000111111111111110000",--28702
"001001111100000000011111111111101111",--28703
"001011111100000001011111111111101110",--28704
"001001111100000000101111111111101101",--28705
"001011111100000001101111111111101100",--28706
"101110010001111000000010100000000000",--28707
"101110001111111000000010000000000000",--28708
"101110000001111000000001100000000000",--28709
"001001111100000111111111111111101011",--28710
"101001111100010111100000000000010110",--28711
"000111000000000000000000001101001100",--28712
"101001111100000111100000000000010110",--28713
"001101111100000111111111111111101011",--28714
"111110000110000000010001100000000000",--28715
"111110000110011000000001100000000000",--28716
"001111111100000001001111111111101100",--28717
"111110001000001000110001100000000000",--28718
"001101111100000000011111111111101101",--28719
"010100000011000000000000000000000100",--28720
"101111001001110001000011111111001001",--28721
"101111001001100001000000111111011010",--28722
"111110001000010000110001100000000000",--28723
"000101000000000000000111000000111001",--28724
"011000000011000000000000000000000011",--28725
"101111001001110001001011111111001001",--28726
"101111001001100001000000111111011010",--28727
"111110001000010000110001100000000000",--28728
"001111111100000001101111111111111101",--28729
"111110000110001001100001100000000000",--28730
"111110000110001000110010000000000000",--28731
"101111000001110001010100000011100000",--28732
"101111001111110001110011110111100011",--28733
"101111001111100001111000111000111001",--28734
"111110001000001001110011100000000000",--28735
"101111000001110010000100000010100000",--28736
"111110001010010001110010100000000000",--28737
"111110001010011000000010100000000000",--28738
"111110001000001001010010100000000000",--28739
"101111000001110001110100000001000000",--28740
"111110010000010001010010100000000000",--28741
"111110001010011000000010100000000000",--28742
"111110001000001001010010100000000000",--28743
"111110001110010001010010100000000000",--28744
"111110001010011000000010100000000000",--28745
"111110001000001001010010000000000000",--28746
"111110001000010000010010000000000010",--28747
"111110001000011000000010000000000000",--28748
"111110000110001001000001100000000000",--28749
"001111111100000001001111111111101110",--28750
"111110000110001001000010000000000000",--28751
"001111111100000000111111111111110000",--28752
"001111111100000001011111111111110010",--28753
"001101111100000000011111111111101111",--28754
"001101111100000000101111111111111110",--28755
"001101111100000000111111111111110100",--28756
"001001111100000111111111111111101011",--28757
"101001111100010111100000000000010110",--28758
"000111000000000000000110110001101000",--28759
"101001111100000111100000000000010110",--28760
"001101111100000111111111111111101011",--28761
"001101111100000000010000000000000000",--28762
"101001000010010000010000000000000001",--28763
"010111000010000000001111100000000000",--28764
"001101111100000000101111111111111110",--28765
"101001000100000000100000000000000001",--28766
"010111000101000001000000000000000001",--28767
"101001000100010000100000000000000101",--28768
"101010000011101000000001100000000000",--28769
"101111001001110001000011111001001100",--28770
"101111001001100001001100110011001101",--28771
"111110000110001001000001100000000000",--28772
"101111001001110001000011111101100110",--28773
"101111001001100001000110011001100110",--28774
"111110000110010001000001100000000000",--28775
"101111001001110001000011111010100001",--28776
"101111001001100001001110100010011001",--28777
"101111001011110001010011111010100001",--28778
"101111001011100001011110100010011000",--28779
"101111001101110001100011110111001100",--28780
"101111001101100001101100110011000101",--28781
"101111010001110010000011110100000101",--28782
"101111010001100010000001001001010001",--28783
"001001111100000000011111111111101011",--28784
"001001111100000000101111111111101010",--28785
"001011111100000001001111111111101001",--28786
"001011111100000000111111111111101000",--28787
"001011111100000001011111111111100111",--28788
"101110010001111000000010100000000000",--28789
"101110001101111000000010000000000000",--28790
"101110000001111000000001100000000000",--28791
"001001111100000111111111111111100110",--28792
"101001111100010111100000000000011011",--28793
"000111000000000000000000001101001100",--28794
"101001111100000111100000000000011011",--28795
"001101111100000111111111111111100110",--28796
"111110000110000000010001100000000000",--28797
"111110000110011000000001100000000000",--28798
"001111111100000001001111111111100111",--28799
"111110001000001000110001100000000000",--28800
"101111001001110001000011111111001001",--28801
"101111001001100001000000111111011010",--28802
"111110001000010000110001100000000000",--28803
"001111111100000001001111111111101000",--28804
"111110000110001001000001100000000000",--28805
"111110000110001000110010100000000000",--28806
"101111000001110001100100000011100000",--28807
"101111001111110001110011110111100011",--28808
"101111001111100001111000111000111001",--28809
"111110001010001001110011100000000000",--28810
"101111000001110010000100000010100000",--28811
"111110001100010001110011000000000000",--28812
"111110001100011000000011000000000000",--28813
"111110001010001001100011000000000000",--28814
"101111000001110001110100000001000000",--28815
"111110010000010001100011000000000000",--28816
"111110001100011000000011000000000000",--28817
"111110001010001001100011000000000000",--28818
"111110001110010001100011000000000000",--28819
"111110001100011000000011000000000000",--28820
"111110001010001001100010100000000000",--28821
"111110001010010000010010100000000010",--28822
"111110001010011000000010100000000000",--28823
"111110000110001001010001100000000000",--28824
"001111111100000001011111111111101001",--28825
"111110000110001001010001100000000000",--28826
"101001000000000000010000000000000001",--28827
"111110000110001000110010100000000000",--28828
"101111001101110001100011110111001100",--28829
"101111001101100001101100110011001101",--28830
"111110001010000001100010100000000000",--28831
"111110001010100000000010100000000000",--28832
"111110001010011000000011000000000000",--28833
"010110001101000000010000000000000010",--28834
"101001000000000000100000000000000001",--28835
"000101000000000000000111000010101010",--28836
"011010001101000000100000000000000010",--28837
"101001000000000000101111111111111111",--28838
"000101000000000000000111000010101010",--28839
"101000000001111000000001000000000000",--28840
"000101000000000000000111000010101011",--28841
"111110001100011000000011000000000000",--28842
"111110001100001001100011100000000000",--28843
"101111000001110010000100001011110010",--28844
"111110010000001001110100000000000000",--28845
"101111010011110010010011110100110010",--28846
"101111010011100010010001011001000011",--28847
"111110010000001010010100000000000000",--28848
"101111000001110010010100001011001000",--28849
"111110010010001001110100100000000000",--28850
"101111000001110010100100000110101000",--28851
"111110010100000010000100000000000000",--28852
"111110010000011000000100000000000000",--28853
"111110010010001010000100000000000000",--28854
"101111000001110010010100001010100010",--28855
"111110010010001001110100100000000000",--28856
"101111000001110010100100000110011000",--28857
"111110010100000010000100000000000000",--28858
"111110010000011000000100000000000000",--28859
"111110010010001010000100000000000000",--28860
"101111000001110010010100001010000000",--28861
"111110010010001001110100100000000000",--28862
"101111000001110010100100000110001000",--28863
"111110010100000010000100000000000000",--28864
"111110010000011000000100000000000000",--28865
"111110010010001010000100000000000000",--28866
"101111000001110010010100001001000100",--28867
"111110010010001001110100100000000000",--28868
"101111000001110010100100000101110000",--28869
"111110010100000010000100000000000000",--28870
"111110010000011000000100000000000000",--28871
"111110010010001010000100000000000000",--28872
"101111000001110010010100001000010000",--28873
"111110010010001001110100100000000000",--28874
"101111000001110010100100000101010000",--28875
"111110010100000010000100000000000000",--28876
"111110010000011000000100000000000000",--28877
"111110010010001010000100000000000000",--28878
"101111000001110010010100000111001000",--28879
"111110010010001001110100100000000000",--28880
"101111000001110010100100000100110000",--28881
"111110010100000010000100000000000000",--28882
"111110010000011000000100000000000000",--28883
"111110010010001010000100000000000000",--28884
"101111000001110010010100000110000000",--28885
"111110010010001001110100100000000000",--28886
"101111000001110010100100000100010000",--28887
"111110010100000010000100000000000000",--28888
"111110010000011000000100000000000000",--28889
"111110010010001010000100000000000000",--28890
"101111000001110010010100000100010000",--28891
"111110010010001001110100100000000000",--28892
"101111000001110010100100000011100000",--28893
"111110010100000010000100000000000000",--28894
"111110010000011000000100000000000000",--28895
"111110010010001010000100000000000000",--28896
"101111000001110010010100000010000000",--28897
"111110010010001001110100100000000000",--28898
"101111000001110010100100000010100000",--28899
"111110010100000010000100000000000000",--28900
"111110010000011000000100000000000000",--28901
"111110010010001010000100000000000000",--28902
"101111000001110010100100000001000000",--28903
"111110010100000010000100000000000000",--28904
"111110010000011000000100000000000000",--28905
"111110001110001010000100000000000000",--28906
"001011111100000000111111111111100110",--28907
"001001111100000000011111111111100101",--28908
"001011111100000001011111111111100100",--28909
"001001111100000000101111111111100011",--28910
"001011111100000001101111111111100010",--28911
"101110010001111000000010100000000000",--28912
"101110001111111000000010000000000000",--28913
"101110000001111000000001100000000000",--28914
"001001111100000111111111111111100001",--28915
"101001111100010111100000000000100000",--28916
"000111000000000000000000001101001100",--28917
"101001111100000111100000000000100000",--28918
"001101111100000111111111111111100001",--28919
"111110000110000000010001100000000000",--28920
"111110000110011000000001100000000000",--28921
"001111111100000001001111111111100010",--28922
"111110001000001000110001100000000000",--28923
"001101111100000000011111111111100011",--28924
"010100000011000000000000000000000100",--28925
"101111001001110001000011111111001001",--28926
"101111001001100001000000111111011010",--28927
"111110001000010000110001100000000000",--28928
"000101000000000000000111000100000110",--28929
"011000000011000000000000000000000011",--28930
"101111001001110001001011111111001001",--28931
"101111001001100001000000111111011010",--28932
"111110001000010000110001100000000000",--28933
"001111111100000001101111111111111101",--28934
"111110000110001001100001100000000000",--28935
"111110000110001000110010000000000000",--28936
"101111000001110001010100000011100000",--28937
"101111001111110001110011110111100011",--28938
"101111001111100001111000111000111001",--28939
"111110001000001001110011100000000000",--28940
"101111000001110010000100000010100000",--28941
"111110001010010001110010100000000000",--28942
"111110001010011000000010100000000000",--28943
"111110001000001001010010100000000000",--28944
"101111000001110001110100000001000000",--28945
"111110010000010001010010100000000000",--28946
"111110001010011000000010100000000000",--28947
"111110001000001001010010100000000000",--28948
"111110001110010001010010100000000000",--28949
"111110001010011000000010100000000000",--28950
"111110001000001001010010000000000000",--28951
"111110001000010000010010000000000010",--28952
"111110001000011000000010000000000000",--28953
"111110000110001001000001100000000000",--28954
"001111111100000001001111111111100100",--28955
"111110000110001001000010000000000000",--28956
"001111111100000000111111111111100110",--28957
"001111111100000001011111111111101000",--28958
"001101111100000000011111111111100101",--28959
"001101111100000000101111111111101010",--28960
"001101111100000000111111111111111111",--28961
"001001111100000111111111111111100001",--28962
"101001111100010111100000000000100000",--28963
"000111000000000000000110110001101000",--28964
"101001111100000111100000000000100000",--28965
"001101111100000111111111111111100001",--28966
"001101111100000000011111111111111111",--28967
"101001000010000000100000000000000010",--28968
"001101111100000000111111111111101011",--28969
"101010000111101000000001100000000000",--28970
"101111001001110001000011111001001100",--28971
"101111001001100001001100110011001101",--28972
"111110000110001001000001100000000000",--28973
"101111001001110001000011110111001100",--28974
"101111001001100001001100110011001101",--28975
"111110000110000001000001100000000000",--28976
"101111001001110001000011111010100001",--28977
"101111001001100001001110100010011001",--28978
"101111001011110001010011111010100001",--28979
"101111001011100001011110100010011000",--28980
"101111001101110001100011110111001100",--28981
"101111001101100001101100110011000101",--28982
"101111010001110010000011110100000101",--28983
"101111010001100010000001001001010001",--28984
"001001111100000000101111111111100001",--28985
"001011111100000001001111111111100000",--28986
"001011111100000000111111111111011111",--28987
"001011111100000001011111111111011110",--28988
"101110010001111000000010100000000000",--28989
"101110001101111000000010000000000000",--28990
"101110000001111000000001100000000000",--28991
"001001111100000111111111111111011101",--28992
"101001111100010111100000000000100100",--28993
"000111000000000000000000001101001100",--28994
"101001111100000111100000000000100100",--28995
"001101111100000111111111111111011101",--28996
"111110000110000000010001100000000000",--28997
"111110000110011000000001100000000000",--28998
"001111111100000001001111111111011110",--28999
"111110001000001000110001100000000000",--29000
"101111001001110001000011111111001001",--29001
"101111001001100001000000111111011010",--29002
"111110001000010000110001100000000000",--29003
"001111111100000001001111111111011111",--29004
"111110000110001001000001100000000000",--29005
"111110000110001000110010100000000000",--29006
"101111000001110001100100000011100000",--29007
"101111001111110001110011110111100011",--29008
"101111001111100001111000111000111001",--29009
"111110001010001001110011100000000000",--29010
"101111000001110010000100000010100000",--29011
"111110001100010001110011000000000000",--29012
"111110001100011000000011000000000000",--29013
"111110001010001001100011000000000000",--29014
"101111000001110001110100000001000000",--29015
"111110010000010001100011000000000000",--29016
"111110001100011000000011000000000000",--29017
"111110001010001001100011000000000000",--29018
"111110001110010001100011000000000000",--29019
"111110001100011000000011000000000000",--29020
"111110001010001001100010100000000000",--29021
"111110001010010000010010100000000010",--29022
"111110001010011000000010100000000000",--29023
"111110000110001001010001100000000000",--29024
"001111111100000001011111111111100000",--29025
"111110000110001001010001100000000000",--29026
"101001000000000000010000000000000001",--29027
"111110000110001000110010100000000000",--29028
"101111001101110001100011110111001100",--29029
"101111001101100001101100110011001101",--29030
"111110001010000001100010100000000000",--29031
"111110001010100000000010100000000000",--29032
"111110001010011000000011000000000000",--29033
"010110001101000000010000000000000010",--29034
"101001000000000000100000000000000001",--29035
"000101000000000000000111000101110010",--29036
"011010001101000000100000000000000010",--29037
"101001000000000000101111111111111111",--29038
"000101000000000000000111000101110010",--29039
"101000000001111000000001000000000000",--29040
"000101000000000000000111000101110011",--29041
"111110001100011000000011000000000000",--29042
"111110001100001001100011100000000000",--29043
"101111000001110010000100001011110010",--29044
"111110010000001001110100000000000000",--29045
"101111010011110010010011110100110010",--29046
"101111010011100010010001011001000011",--29047
"111110010000001010010100000000000000",--29048
"101111000001110010010100001011001000",--29049
"111110010010001001110100100000000000",--29050
"101111000001110010100100000110101000",--29051
"111110010100000010000100000000000000",--29052
"111110010000011000000100000000000000",--29053
"111110010010001010000100000000000000",--29054
"101111000001110010010100001010100010",--29055
"111110010010001001110100100000000000",--29056
"101111000001110010100100000110011000",--29057
"111110010100000010000100000000000000",--29058
"111110010000011000000100000000000000",--29059
"111110010010001010000100000000000000",--29060
"101111000001110010010100001010000000",--29061
"111110010010001001110100100000000000",--29062
"101111000001110010100100000110001000",--29063
"111110010100000010000100000000000000",--29064
"111110010000011000000100000000000000",--29065
"111110010010001010000100000000000000",--29066
"101111000001110010010100001001000100",--29067
"111110010010001001110100100000000000",--29068
"101111000001110010100100000101110000",--29069
"111110010100000010000100000000000000",--29070
"111110010000011000000100000000000000",--29071
"111110010010001010000100000000000000",--29072
"101111000001110010010100001000010000",--29073
"111110010010001001110100100000000000",--29074
"101111000001110010100100000101010000",--29075
"111110010100000010000100000000000000",--29076
"111110010000011000000100000000000000",--29077
"111110010010001010000100000000000000",--29078
"101111000001110010010100000111001000",--29079
"111110010010001001110100100000000000",--29080
"101111000001110010100100000100110000",--29081
"111110010100000010000100000000000000",--29082
"111110010000011000000100000000000000",--29083
"111110010010001010000100000000000000",--29084
"101111000001110010010100000110000000",--29085
"111110010010001001110100100000000000",--29086
"101111000001110010100100000100010000",--29087
"111110010100000010000100000000000000",--29088
"111110010000011000000100000000000000",--29089
"111110010010001010000100000000000000",--29090
"101111000001110010010100000100010000",--29091
"111110010010001001110100100000000000",--29092
"101111000001110010100100000011100000",--29093
"111110010100000010000100000000000000",--29094
"111110010000011000000100000000000000",--29095
"111110010010001010000100000000000000",--29096
"101111000001110010010100000010000000",--29097
"111110010010001001110100100000000000",--29098
"101111000001110010100100000010100000",--29099
"111110010100000010000100000000000000",--29100
"111110010000011000000100000000000000",--29101
"111110010010001010000100000000000000",--29102
"101111000001110010100100000001000000",--29103
"111110010100000010000100000000000000",--29104
"111110010000011000000100000000000000",--29105
"111110001110001010000100000000000000",--29106
"001011111100000000111111111111011101",--29107
"001001111100000000011111111111011100",--29108
"001011111100000001011111111111011011",--29109
"001001111100000000101111111111011010",--29110
"001011111100000001101111111111011001",--29111
"101110010001111000000010100000000000",--29112
"101110001111111000000010000000000000",--29113
"101110000001111000000001100000000000",--29114
"001001111100000111111111111111011000",--29115
"101001111100010111100000000000101001",--29116
"000111000000000000000000001101001100",--29117
"101001111100000111100000000000101001",--29118
"001101111100000111111111111111011000",--29119
"111110000110000000010001100000000000",--29120
"111110000110011000000001100000000000",--29121
"001111111100000001001111111111011001",--29122
"111110001000001000110001100000000000",--29123
"001101111100000000011111111111011010",--29124
"010100000011000000000000000000000100",--29125
"101111001001110001000011111111001001",--29126
"101111001001100001000000111111011010",--29127
"111110001000010000110001100000000000",--29128
"000101000000000000000111000111001110",--29129
"011000000011000000000000000000000011",--29130
"101111001001110001001011111111001001",--29131
"101111001001100001000000111111011010",--29132
"111110001000010000110001100000000000",--29133
"001111111100000001101111111111111101",--29134
"111110000110001001100001100000000000",--29135
"111110000110001000110010000000000000",--29136
"101111000001110001010100000011100000",--29137
"101111001111110001110011110111100011",--29138
"101111001111100001111000111000111001",--29139
"111110001000001001110011100000000000",--29140
"101111000001110010000100000010100000",--29141
"111110001010010001110010100000000000",--29142
"111110001010011000000010100000000000",--29143
"111110001000001001010010100000000000",--29144
"101111000001110001110100000001000000",--29145
"111110010000010001010010100000000000",--29146
"111110001010011000000010100000000000",--29147
"111110001000001001010010100000000000",--29148
"111110001110010001010010100000000000",--29149
"111110001010011000000010100000000000",--29150
"111110001000001001010010000000000000",--29151
"111110001000010000010010000000000010",--29152
"111110001000011000000010000000000000",--29153
"111110000110001001000001100000000000",--29154
"001111111100000001001111111111011011",--29155
"111110000110001001000010000000000000",--29156
"001111111100000000111111111111011101",--29157
"001111111100000001011111111111011111",--29158
"001101111100000000011111111111011100",--29159
"001101111100000000101111111111101010",--29160
"001101111100000000111111111111100001",--29161
"001001111100000111111111111111011000",--29162
"101001111100010111100000000000101001",--29163
"000111000000000000000110110001101000",--29164
"101001111100000111100000000000101001",--29165
"001101111100000111111111111111011000",--29166
"001101111100000000011111111111101011",--29167
"101001000010010000010000000000000001",--29168
"010111000010000000001111100000000000",--29169
"001101111100000000101111111111101010",--29170
"101001000100000000100000000000000001",--29171
"010111000101000001000000000000000001",--29172
"101001000100010000100000000000000101",--29173
"101010000011101000000001100000000000",--29174
"101111001001110001000011111001001100",--29175
"101111001001100001001100110011001101",--29176
"111110000110001001000001100000000000",--29177
"101111001001110001000011111101100110",--29178
"101111001001100001000110011001100110",--29179
"111110000110010001000010100000000000",--29180
"101110000001111000000001100000000000",--29181
"101110000001111000000010000000000000",--29182
"001111111100000001101111111111111101",--29183
"001101111100000000111111111111111111",--29184
"001001111100000000101111111111011000",--29185
"001001111100000000011111111111010111",--29186
"101000000001111000000000100000000000",--29187
"001001111100000111111111111111010110",--29188
"101001111100010111100000000000101011",--29189
"000111000000000000000110110001101000",--29190
"101001111100000111100000000000101011",--29191
"001101111100000000011111111111010111",--29192
"101010000011101000000001100000000000",--29193
"101111001001110001000011111001001100",--29194
"101111001001100001001100110011001101",--29195
"111110000110001001000001100000000000",--29196
"101111001001110001000011110111001100",--29197
"101111001001100001001100110011001101",--29198
"111110000110000001000010100000000000",--29199
"101110000001111000000001100000000000",--29200
"101110000001111000000010000000000000",--29201
"001101111100000000111111111111111111",--29202
"101001000110000000110000000000000010",--29203
"001111111100000001101111111111111101",--29204
"001101111100000000101111111111011000",--29205
"101000000001111000000000100000000000",--29206
"101001111100010111100000000000101011",--29207
"000111000000000000000110110001101000",--29208
"101001111100000111100000000000101011",--29209
"001101111100000111111111111111010110",--29210
"001101111100000000011111111111010111",--29211
"101001000010010000010000000000000001",--29212
"010111000010000000001111100000000000",--29213
"001101111100000000101111111111011000",--29214
"101001000100000000100000000000000001",--29215
"010111000101000001000000000000000001",--29216
"101001000100010000100000000000000101",--29217
"101010000011101000000001100000000000",--29218
"101111001001110001000011111001001100",--29219
"101111001001100001001100110011001101",--29220
"111110000110001001000001100000000000",--29221
"101111001001110001000011111101100110",--29222
"101111001001100001000110011001100110",--29223
"111110000110010001000010100000000000",--29224
"101110000001111000000001100000000000",--29225
"101110000001111000000010000000000000",--29226
"001111111100000001101111111111111101",--29227
"001101111100000000111111111111111111",--29228
"001001111100000000101111111111010110",--29229
"001001111100000000011111111111010101",--29230
"101000000001111000000000100000000000",--29231
"001001111100000111111111111111010100",--29232
"101001111100010111100000000000101101",--29233
"000111000000000000000110110001101000",--29234
"101001111100000111100000000000101101",--29235
"001101111100000000011111111111010101",--29236
"101010000011101000000001100000000000",--29237
"101111001001110001000011111001001100",--29238
"101111001001100001001100110011001101",--29239
"111110000110001001000001100000000000",--29240
"101111001001110001000011110111001100",--29241
"101111001001100001001100110011001101",--29242
"111110000110000001000010100000000000",--29243
"101110000001111000000001100000000000",--29244
"101110000001111000000010000000000000",--29245
"001101111100000000111111111111111111",--29246
"101001000110000000110000000000000010",--29247
"001111111100000001101111111111111101",--29248
"001101111100000000101111111111010110",--29249
"101000000001111000000000100000000000",--29250
"101001111100010111100000000000101101",--29251
"000111000000000000000110110001101000",--29252
"101001111100000111100000000000101101",--29253
"001101111100000111111111111111010100",--29254
"001101111100000000011111111111010101",--29255
"101001000010010000010000000000000001",--29256
"001101111100000000101111111111010110",--29257
"101001000100000000100000000000000001",--29258
"010111000101000001000000000000000001",--29259
"101001000100010000100000000000000101",--29260
"001111111100000000111111111111111101",--29261
"001101111100000000111111111111111111",--29262
"010111000010000000001111100000000000",--29263
"000101000000000000000110111011001010",--29264
"010111000010000000001111100000000000",--29265
"101001000000000001000000000000000100",--29266
"101010000011101000000001100000000000",--29267
"101111001001110001000011111001001100",--29268
"101111001001100001001100110011001101",--29269
"111110000110001001000001100000000000",--29270
"101111001001110001000011111101100110",--29271
"101111001001100001000110011001100110",--29272
"111110000110010001000001100000000000",--29273
"101010001001101000000010000000000000",--29274
"101111001011110001010011111001001100",--29275
"101111001011100001011100110011001101",--29276
"111110001000001001010010000000000000",--29277
"101111001011110001010011111101100110",--29278
"101111001011100001010110011001100110",--29279
"111110001000010001010010000000000000",--29280
"101111001011110001010011111010100001",--29281
"101111001011100001011110100010011001",--29282
"101111001101110001100011111010100001",--29283
"101111001101100001101110100010011000",--29284
"101111001111110001110011110111001100",--29285
"101111001111100001111100110011000101",--29286
"101111010011110010010011110100000101",--29287
"101111010011100010010001001001010001",--29288
"001001111100000000010000000000000000",--29289
"001001111100000001001111111111111111",--29290
"001001111100000000111111111111111110",--29291
"001001111100000000101111111111111101",--29292
"001011111100000000111111111111111100",--29293
"001011111100000001011111111111111011",--29294
"001011111100000001001111111111111010",--29295
"001011111100000001101111111111111001",--29296
"101110010011111000000010100000000000",--29297
"101110001111111000000010000000000000",--29298
"101110000001111000000001100000000000",--29299
"001001111100000111111111111111111000",--29300
"101001111100010111100000000000001001",--29301
"000111000000000000000000001101001100",--29302
"101001111100000111100000000000001001",--29303
"001101111100000111111111111111111000",--29304
"111110000110000000010001100000000000",--29305
"111110000110011000000001100000000000",--29306
"001111111100000001001111111111111001",--29307
"111110001000001000110001100000000000",--29308
"101111001001110001000011111111001001",--29309
"101111001001100001000000111111011010",--29310
"111110001000010000110001100000000000",--29311
"001111111100000001001111111111111010",--29312
"111110000110001001000001100000000000",--29313
"111110000110001000110010100000000000",--29314
"101111000001110001100100000011100000",--29315
"101111001111110001110011110111100011",--29316
"101111001111100001111000111000111001",--29317
"111110001010001001110011100000000000",--29318
"101111000001110010000100000010100000",--29319
"111110001100010001110011000000000000",--29320
"111110001100011000000011000000000000",--29321
"111110001010001001100011000000000000",--29322
"101111000001110001110100000001000000",--29323
"111110010000010001100011000000000000",--29324
"111110001100011000000011000000000000",--29325
"111110001010001001100011000000000000",--29326
"111110001110010001100011000000000000",--29327
"111110001100011000000011000000000000",--29328
"111110001010001001100010100000000000",--29329
"111110001010010000010010100000000010",--29330
"111110001010011000000010100000000000",--29331
"111110000110001001010001100000000000",--29332
"001111111100000001011111111111111011",--29333
"111110000110001001010001100000000000",--29334
"101001000000000000010000000000000001",--29335
"111110000110001000110010100000000000",--29336
"101111001101110001100011110111001100",--29337
"101111001101100001101100110011001101",--29338
"111110001010000001100010100000000000",--29339
"111110001010100000000010100000000000",--29340
"111110001010011000000011000000000000",--29341
"010110001101000000010000000000000010",--29342
"101001000000000000100000000000000001",--29343
"000101000000000000000111001010100110",--29344
"011010001101000000100000000000000010",--29345
"101001000000000000101111111111111111",--29346
"000101000000000000000111001010100110",--29347
"101000000001111000000001000000000000",--29348
"000101000000000000000111001010100111",--29349
"111110001100011000000011000000000000",--29350
"111110001100001001100011100000000000",--29351
"101111000001110010000100001011110010",--29352
"111110010000001001110100000000000000",--29353
"101111010011110010010011110100110010",--29354
"101111010011100010010001011001000011",--29355
"111110010000001010010100000000000000",--29356
"101111000001110010010100001011001000",--29357
"111110010010001001110100100000000000",--29358
"101111000001110010100100000110101000",--29359
"111110010100000010000100000000000000",--29360
"111110010000011000000100000000000000",--29361
"111110010010001010000100000000000000",--29362
"101111000001110010010100001010100010",--29363
"111110010010001001110100100000000000",--29364
"101111000001110010100100000110011000",--29365
"111110010100000010000100000000000000",--29366
"111110010000011000000100000000000000",--29367
"111110010010001010000100000000000000",--29368
"101111000001110010010100001010000000",--29369
"111110010010001001110100100000000000",--29370
"101111000001110010100100000110001000",--29371
"111110010100000010000100000000000000",--29372
"111110010000011000000100000000000000",--29373
"111110010010001010000100000000000000",--29374
"101111000001110010010100001001000100",--29375
"111110010010001001110100100000000000",--29376
"101111000001110010100100000101110000",--29377
"111110010100000010000100000000000000",--29378
"111110010000011000000100000000000000",--29379
"111110010010001010000100000000000000",--29380
"101111000001110010010100001000010000",--29381
"111110010010001001110100100000000000",--29382
"101111000001110010100100000101010000",--29383
"111110010100000010000100000000000000",--29384
"111110010000011000000100000000000000",--29385
"111110010010001010000100000000000000",--29386
"101111000001110010010100000111001000",--29387
"111110010010001001110100100000000000",--29388
"101111000001110010100100000100110000",--29389
"111110010100000010000100000000000000",--29390
"111110010000011000000100000000000000",--29391
"111110010010001010000100000000000000",--29392
"101111000001110010010100000110000000",--29393
"111110010010001001110100100000000000",--29394
"101111000001110010100100000100010000",--29395
"111110010100000010000100000000000000",--29396
"111110010000011000000100000000000000",--29397
"111110010010001010000100000000000000",--29398
"101111000001110010010100000100010000",--29399
"111110010010001001110100100000000000",--29400
"101111000001110010100100000011100000",--29401
"111110010100000010000100000000000000",--29402
"111110010000011000000100000000000000",--29403
"111110010010001010000100000000000000",--29404
"101111000001110010010100000010000000",--29405
"111110010010001001110100100000000000",--29406
"101111000001110010100100000010100000",--29407
"111110010100000010000100000000000000",--29408
"111110010000011000000100000000000000",--29409
"111110010010001010000100000000000000",--29410
"101111000001110010100100000001000000",--29411
"111110010100000010000100000000000000",--29412
"111110010000011000000100000000000000",--29413
"111110001110001010000100000000000000",--29414
"001011111100000000111111111111111000",--29415
"001001111100000000011111111111110111",--29416
"001011111100000001011111111111110110",--29417
"001001111100000000101111111111110101",--29418
"001011111100000001101111111111110100",--29419
"101110010001111000000010100000000000",--29420
"101110001111111000000010000000000000",--29421
"101110000001111000000001100000000000",--29422
"001001111100000111111111111111110011",--29423
"101001111100010111100000000000001110",--29424
"000111000000000000000000001101001100",--29425
"101001111100000111100000000000001110",--29426
"001101111100000111111111111111110011",--29427
"111110000110000000010001100000000000",--29428
"111110000110011000000001100000000000",--29429
"001111111100000001001111111111110100",--29430
"111110001000001000110001100000000000",--29431
"001101111100000000011111111111110101",--29432
"010100000011000000000000000000000100",--29433
"101111001001110001000011111111001001",--29434
"101111001001100001000000111111011010",--29435
"111110001000010000110001100000000000",--29436
"000101000000000000000111001100000010",--29437
"011000000011000000000000000000000011",--29438
"101111001001110001001011111111001001",--29439
"101111001001100001000000111111011010",--29440
"111110001000010000110001100000000000",--29441
"001111111100000001101111111111111100",--29442
"111110000110001001100001100000000000",--29443
"111110000110001000110010000000000000",--29444
"101111000001110001010100000011100000",--29445
"101111001111110001110011110111100011",--29446
"101111001111100001111000111000111001",--29447
"111110001000001001110011100000000000",--29448
"101111000001110010000100000010100000",--29449
"111110001010010001110010100000000000",--29450
"111110001010011000000010100000000000",--29451
"111110001000001001010010100000000000",--29452
"101111000001110001110100000001000000",--29453
"111110010000010001010010100000000000",--29454
"111110001010011000000010100000000000",--29455
"111110001000001001010010100000000000",--29456
"111110001110010001010010100000000000",--29457
"111110001010011000000010100000000000",--29458
"111110001000001001010010000000000000",--29459
"111110001000010000010010000000000010",--29460
"111110001000011000000010000000000000",--29461
"111110000110001001000001100000000000",--29462
"001111111100000001001111111111110110",--29463
"111110000110001001000010000000000000",--29464
"001111111100000000111111111111111000",--29465
"001111111100000001011111111111111010",--29466
"001101111100000000011111111111110111",--29467
"001101111100000000101111111111111101",--29468
"001101111100000000111111111111111110",--29469
"001001111100000111111111111111110011",--29470
"101001111100010111100000000000001110",--29471
"000111000000000000000110110001101000",--29472
"101001111100000111100000000000001110",--29473
"001101111100000111111111111111110011",--29474
"001101111100000000011111111111111110",--29475
"101001000010000000100000000000000010",--29476
"001101111100000000111111111111111111",--29477
"101010000111101000000001100000000000",--29478
"101111001001110001000011111001001100",--29479
"101111001001100001001100110011001101",--29480
"111110000110001001000001100000000000",--29481
"101111001001110001000011110111001100",--29482
"101111001001100001001100110011001101",--29483
"111110000110000001000001100000000000",--29484
"101111001001110001000011111010100001",--29485
"101111001001100001001110100010011001",--29486
"101111001011110001010011111010100001",--29487
"101111001011100001011110100010011000",--29488
"101111001101110001100011110111001100",--29489
"101111001101100001101100110011000101",--29490
"101111010001110010000011110100000101",--29491
"101111010001100010000001001001010001",--29492
"001001111100000000101111111111110011",--29493
"001011111100000001001111111111110010",--29494
"001011111100000000111111111111110001",--29495
"001011111100000001011111111111110000",--29496
"101110010001111000000010100000000000",--29497
"101110001101111000000010000000000000",--29498
"101110000001111000000001100000000000",--29499
"001001111100000111111111111111101111",--29500
"101001111100010111100000000000010010",--29501
"000111000000000000000000001101001100",--29502
"101001111100000111100000000000010010",--29503
"001101111100000111111111111111101111",--29504
"111110000110000000010001100000000000",--29505
"111110000110011000000001100000000000",--29506
"001111111100000001001111111111110000",--29507
"111110001000001000110001100000000000",--29508
"101111001001110001000011111111001001",--29509
"101111001001100001000000111111011010",--29510
"111110001000010000110001100000000000",--29511
"001111111100000001001111111111110001",--29512
"111110000110001001000001100000000000",--29513
"111110000110001000110010100000000000",--29514
"101111000001110001100100000011100000",--29515
"101111001111110001110011110111100011",--29516
"101111001111100001111000111000111001",--29517
"111110001010001001110011100000000000",--29518
"101111000001110010000100000010100000",--29519
"111110001100010001110011000000000000",--29520
"111110001100011000000011000000000000",--29521
"111110001010001001100011000000000000",--29522
"101111000001110001110100000001000000",--29523
"111110010000010001100011000000000000",--29524
"111110001100011000000011000000000000",--29525
"111110001010001001100011000000000000",--29526
"111110001110010001100011000000000000",--29527
"111110001100011000000011000000000000",--29528
"111110001010001001100010100000000000",--29529
"111110001010010000010010100000000010",--29530
"111110001010011000000010100000000000",--29531
"111110000110001001010001100000000000",--29532
"001111111100000001011111111111110010",--29533
"111110000110001001010001100000000000",--29534
"101001000000000000010000000000000001",--29535
"111110000110001000110010100000000000",--29536
"101111001101110001100011110111001100",--29537
"101111001101100001101100110011001101",--29538
"111110001010000001100010100000000000",--29539
"111110001010100000000010100000000000",--29540
"111110001010011000000011000000000000",--29541
"010110001101000000010000000000000010",--29542
"101001000000000000100000000000000001",--29543
"000101000000000000000111001101101110",--29544
"011010001101000000100000000000000010",--29545
"101001000000000000101111111111111111",--29546
"000101000000000000000111001101101110",--29547
"101000000001111000000001000000000000",--29548
"000101000000000000000111001101101111",--29549
"111110001100011000000011000000000000",--29550
"111110001100001001100011100000000000",--29551
"101111000001110010000100001011110010",--29552
"111110010000001001110100000000000000",--29553
"101111010011110010010011110100110010",--29554
"101111010011100010010001011001000011",--29555
"111110010000001010010100000000000000",--29556
"101111000001110010010100001011001000",--29557
"111110010010001001110100100000000000",--29558
"101111000001110010100100000110101000",--29559
"111110010100000010000100000000000000",--29560
"111110010000011000000100000000000000",--29561
"111110010010001010000100000000000000",--29562
"101111000001110010010100001010100010",--29563
"111110010010001001110100100000000000",--29564
"101111000001110010100100000110011000",--29565
"111110010100000010000100000000000000",--29566
"111110010000011000000100000000000000",--29567
"111110010010001010000100000000000000",--29568
"101111000001110010010100001010000000",--29569
"111110010010001001110100100000000000",--29570
"101111000001110010100100000110001000",--29571
"111110010100000010000100000000000000",--29572
"111110010000011000000100000000000000",--29573
"111110010010001010000100000000000000",--29574
"101111000001110010010100001001000100",--29575
"111110010010001001110100100000000000",--29576
"101111000001110010100100000101110000",--29577
"111110010100000010000100000000000000",--29578
"111110010000011000000100000000000000",--29579
"111110010010001010000100000000000000",--29580
"101111000001110010010100001000010000",--29581
"111110010010001001110100100000000000",--29582
"101111000001110010100100000101010000",--29583
"111110010100000010000100000000000000",--29584
"111110010000011000000100000000000000",--29585
"111110010010001010000100000000000000",--29586
"101111000001110010010100000111001000",--29587
"111110010010001001110100100000000000",--29588
"101111000001110010100100000100110000",--29589
"111110010100000010000100000000000000",--29590
"111110010000011000000100000000000000",--29591
"111110010010001010000100000000000000",--29592
"101111000001110010010100000110000000",--29593
"111110010010001001110100100000000000",--29594
"101111000001110010100100000100010000",--29595
"111110010100000010000100000000000000",--29596
"111110010000011000000100000000000000",--29597
"111110010010001010000100000000000000",--29598
"101111000001110010010100000100010000",--29599
"111110010010001001110100100000000000",--29600
"101111000001110010100100000011100000",--29601
"111110010100000010000100000000000000",--29602
"111110010000011000000100000000000000",--29603
"111110010010001010000100000000000000",--29604
"101111000001110010010100000010000000",--29605
"111110010010001001110100100000000000",--29606
"101111000001110010100100000010100000",--29607
"111110010100000010000100000000000000",--29608
"111110010000011000000100000000000000",--29609
"111110010010001010000100000000000000",--29610
"101111000001110010100100000001000000",--29611
"111110010100000010000100000000000000",--29612
"111110010000011000000100000000000000",--29613
"111110001110001010000100000000000000",--29614
"001011111100000000111111111111101111",--29615
"001001111100000000011111111111101110",--29616
"001011111100000001011111111111101101",--29617
"001001111100000000101111111111101100",--29618
"001011111100000001101111111111101011",--29619
"101110010001111000000010100000000000",--29620
"101110001111111000000010000000000000",--29621
"101110000001111000000001100000000000",--29622
"001001111100000111111111111111101010",--29623
"101001111100010111100000000000010111",--29624
"000111000000000000000000001101001100",--29625
"101001111100000111100000000000010111",--29626
"001101111100000111111111111111101010",--29627
"111110000110000000010001100000000000",--29628
"111110000110011000000001100000000000",--29629
"001111111100000001001111111111101011",--29630
"111110001000001000110001100000000000",--29631
"001101111100000000011111111111101100",--29632
"010100000011000000000000000000000100",--29633
"101111001001110001000011111111001001",--29634
"101111001001100001000000111111011010",--29635
"111110001000010000110001100000000000",--29636
"000101000000000000000111001111001010",--29637
"011000000011000000000000000000000011",--29638
"101111001001110001001011111111001001",--29639
"101111001001100001000000111111011010",--29640
"111110001000010000110001100000000000",--29641
"001111111100000001101111111111111100",--29642
"111110000110001001100001100000000000",--29643
"111110000110001000110010000000000000",--29644
"101111000001110001010100000011100000",--29645
"101111001111110001110011110111100011",--29646
"101111001111100001111000111000111001",--29647
"111110001000001001110011100000000000",--29648
"101111000001110010000100000010100000",--29649
"111110001010010001110010100000000000",--29650
"111110001010011000000010100000000000",--29651
"111110001000001001010010100000000000",--29652
"101111000001110001110100000001000000",--29653
"111110010000010001010010100000000000",--29654
"111110001010011000000010100000000000",--29655
"111110001000001001010010100000000000",--29656
"111110001110010001010010100000000000",--29657
"111110001010011000000010100000000000",--29658
"111110001000001001010010000000000000",--29659
"111110001000010000010010000000000010",--29660
"111110001000011000000010000000000000",--29661
"111110000110001001000001100000000000",--29662
"001111111100000001001111111111101101",--29663
"111110000110001001000010000000000000",--29664
"001111111100000000111111111111101111",--29665
"001111111100000001011111111111110001",--29666
"001101111100000000011111111111101110",--29667
"001101111100000000101111111111111101",--29668
"001101111100000000111111111111110011",--29669
"001001111100000111111111111111101010",--29670
"101001111100010111100000000000010111",--29671
"000111000000000000000110110001101000",--29672
"101001111100000111100000000000010111",--29673
"001101111100000111111111111111101010",--29674
"101001000000000000010000000000000011",--29675
"001101111100000000101111111111111101",--29676
"101001000100000000110000000000000001",--29677
"010111000111000001000000000000000001",--29678
"101001000110010000110000000000000101",--29679
"101010000011101000000001100000000000",--29680
"101111001001110001000011111001001100",--29681
"101111001001100001001100110011001101",--29682
"111110000110001001000001100000000000",--29683
"101111001001110001000011111101100110",--29684
"101111001001100001000110011001100110",--29685
"111110000110010001000010100000000000",--29686
"101110000001111000000001100000000000",--29687
"101110000001111000000010000000000000",--29688
"001111111100000001101111111111111100",--29689
"001101111100000001011111111111111110",--29690
"001001111100000000111111111111101010",--29691
"001001111100000000011111111111101001",--29692
"101000000111111000000001000000000000",--29693
"101000000001111000000000100000000000",--29694
"101000001011111000000001100000000000",--29695
"001001111100000111111111111111101000",--29696
"101001111100010111100000000000011001",--29697
"000111000000000000000110110001101000",--29698
"101001111100000111100000000000011001",--29699
"001101111100000000011111111111101001",--29700
"101010000011101000000001100000000000",--29701
"101111001001110001000011111001001100",--29702
"101111001001100001001100110011001101",--29703
"111110000110001001000001100000000000",--29704
"101111001001110001000011110111001100",--29705
"101111001001100001001100110011001101",--29706
"111110000110000001000010100000000000",--29707
"101000000001111000000000100000000000",--29708
"101110000001111000000001100000000000",--29709
"101110000001111000000010000000000000",--29710
"001101111100000000101111111111111110",--29711
"101001000100000000110000000000000010",--29712
"001111111100000001101111111111111100",--29713
"001101111100000000101111111111101010",--29714
"101001111100010111100000000000011001",--29715
"000111000000000000000110110001101000",--29716
"101001111100000111100000000000011001",--29717
"001101111100000111111111111111101000",--29718
"101001000000000000010000000000000010",--29719
"001101111100000000101111111111101010",--29720
"101001000100000000100000000000000001",--29721
"010111000101000001000000000000000001",--29722
"101001000100010000100000000000000101",--29723
"101010000011101000000001100000000000",--29724
"101111001001110001000011111001001100",--29725
"101111001001100001001100110011001101",--29726
"111110000110001001000001100000000000",--29727
"101111001001110001000011111101100110",--29728
"101111001001100001000110011001100110",--29729
"111110000110010001000010100000000000",--29730
"101110000001111000000001100000000000",--29731
"101110000001111000000010000000000000",--29732
"001111111100000001101111111111111100",--29733
"001101111100000000111111111111111110",--29734
"001001111100000000101111111111101000",--29735
"001001111100000000011111111111100111",--29736
"101000000001111000000000100000000000",--29737
"001001111100000111111111111111100110",--29738
"101001111100010111100000000000011011",--29739
"000111000000000000000110110001101000",--29740
"101001111100000111100000000000011011",--29741
"001101111100000000011111111111100111",--29742
"101010000011101000000001100000000000",--29743
"101111001001110001000011111001001100",--29744
"101111001001100001001100110011001101",--29745
"111110000110001001000001100000000000",--29746
"101111001001110001000011110111001100",--29747
"101111001001100001001100110011001101",--29748
"111110000110000001000010100000000000",--29749
"101000000001111000000000100000000000",--29750
"101110000001111000000001100000000000",--29751
"101110000001111000000010000000000000",--29752
"001101111100000000101111111111111110",--29753
"101001000100000000110000000000000010",--29754
"001111111100000001101111111111111100",--29755
"001101111100000000101111111111101000",--29756
"101001111100010111100000000000011011",--29757
"000111000000000000000110110001101000",--29758
"101001111100000111100000000000011011",--29759
"001101111100000111111111111111100110",--29760
"101001000000000000010000000000000001",--29761
"001101111100000000101111111111101000",--29762
"101001000100000000100000000000000001",--29763
"010111000101000001000000000000000001",--29764
"101001000100010000100000000000000101",--29765
"001111111100000000111111111111111100",--29766
"001101111100000000111111111111111110",--29767
"001001111100000111111111111111100110",--29768
"101001111100010111100000000000011011",--29769
"000111000000000000000110111011001001",--29770
"101001111100000111100000000000011011",--29771
"001101111100000111111111111111100110",--29772
"001101111100000000010000000000000000",--29773
"101001000010010000010000000000000001",--29774
"010111000010000000001111100000000000",--29775
"001101111100000000101111111111111101",--29776
"101001000100000000100000000000000010",--29777
"010111000101000001000000000000000001",--29778
"101001000100010000100000000000000101",--29779
"001101111100000000111111111111111110",--29780
"101001000110000000110000000000000100",--29781
"101001000000000001000000000000000100",--29782
"101010000011101000000001100000000000",--29783
"101111001001110001000011111001001100",--29784
"101111001001100001001100110011001101",--29785
"111110000110001001000001100000000000",--29786
"101111001001110001000011111101100110",--29787
"101111001001100001000110011001100110",--29788
"111110000110010001000011000000000000",--29789
"101010001001101000000001100000000000",--29790
"101111001001110001000011111001001100",--29791
"101111001001100001001100110011001101",--29792
"111110000110001001000001100000000000",--29793
"101111001001110001000011111101100110",--29794
"101111001001100001000110011001100110",--29795
"111110000110010001000010100000000000",--29796
"101110000001111000000001100000000000",--29797
"101110000001111000000010000000000000",--29798
"001001111100000000011111111111100110",--29799
"001011111100000001101111111111100101",--29800
"001001111100000000101111111111100100",--29801
"001001111100000000111111111111100011",--29802
"001001111100000001001111111111100010",--29803
"101000000001111000000000100000000000",--29804
"001001111100000111111111111111100001",--29805
"101001111100010111100000000000100000",--29806
"000111000000000000000110110001101000",--29807
"101001111100000111100000000000100000",--29808
"001101111100000000011111111111100010",--29809
"101010000011101000000001100000000000",--29810
"101111001001110001000011111001001100",--29811
"101111001001100001001100110011001101",--29812
"111110000110001001000001100000000000",--29813
"101111001001110001000011110111001100",--29814
"101111001001100001001100110011001101",--29815
"111110000110000001000010100000000000",--29816
"101000000001111000000000100000000000",--29817
"101110000001111000000001100000000000",--29818
"101110000001111000000010000000000000",--29819
"001101111100000000101111111111100011",--29820
"101001000100000000110000000000000010",--29821
"001111111100000001101111111111100101",--29822
"001101111100000000101111111111100100",--29823
"101001111100010111100000000000100000",--29824
"000111000000000000000110110001101000",--29825
"101001111100000111100000000000100000",--29826
"001101111100000111111111111111100001",--29827
"101001000000000000010000000000000011",--29828
"001101111100000000101111111111100100",--29829
"101001000100000000110000000000000001",--29830
"010111000111000001000000000000000001",--29831
"101001000110010000110000000000000101",--29832
"101010000011101000000001100000000000",--29833
"101111001001110001000011111001001100",--29834
"101111001001100001001100110011001101",--29835
"111110000110001001000001100000000000",--29836
"101111001001110001000011111101100110",--29837
"101111001001100001000110011001100110",--29838
"111110000110010001000010100000000000",--29839
"101110000001111000000001100000000000",--29840
"101110000001111000000010000000000000",--29841
"001111111100000001101111111111100101",--29842
"001101111100000001011111111111100011",--29843
"001001111100000000111111111111100001",--29844
"001001111100000000011111111111100000",--29845
"101000000111111000000001000000000000",--29846
"101000000001111000000000100000000000",--29847
"101000001011111000000001100000000000",--29848
"001001111100000111111111111111011111",--29849
"101001111100010111100000000000100010",--29850
"000111000000000000000110110001101000",--29851
"101001111100000111100000000000100010",--29852
"001101111100000000011111111111100000",--29853
"101010000011101000000001100000000000",--29854
"101111001001110001000011111001001100",--29855
"101111001001100001001100110011001101",--29856
"111110000110001001000001100000000000",--29857
"101111001001110001000011110111001100",--29858
"101111001001100001001100110011001101",--29859
"111110000110000001000010100000000000",--29860
"101000000001111000000000100000000000",--29861
"101110000001111000000001100000000000",--29862
"101110000001111000000010000000000000",--29863
"001101111100000000101111111111100011",--29864
"101001000100000000110000000000000010",--29865
"001111111100000001101111111111100101",--29866
"001101111100000000101111111111100001",--29867
"101001111100010111100000000000100010",--29868
"000111000000000000000110110001101000",--29869
"101001111100000111100000000000100010",--29870
"001101111100000111111111111111011111",--29871
"101001000000000000010000000000000010",--29872
"001101111100000000101111111111100001",--29873
"101001000100000000100000000000000001",--29874
"010111000101000001000000000000000001",--29875
"101001000100010000100000000000000101",--29876
"001111111100000000111111111111100101",--29877
"001101111100000000111111111111100011",--29878
"001001111100000111111111111111011111",--29879
"101001111100010111100000000000100010",--29880
"000111000000000000000110111011001001",--29881
"101001111100000111100000000000100010",--29882
"001101111100000111111111111111011111",--29883
"001101111100000000011111111111100110",--29884
"101001000010010000010000000000000001",--29885
"010111000010000000001111100000000000",--29886
"001101111100000000101111111111100100",--29887
"101001000100000000100000000000000010",--29888
"010111000101000001000000000000000001",--29889
"101001000100010000100000000000000101",--29890
"001101111100000000111111111111100011",--29891
"101001000110000000110000000000000100",--29892
"101001000000000001000000000000000100",--29893
"101010000011101000000001100000000000",--29894
"101111001001110001000011111001001100",--29895
"101111001001100001001100110011001101",--29896
"111110000110001001000001100000000000",--29897
"101111001001110001000011111101100110",--29898
"101111001001100001000110011001100110",--29899
"111110000110010001000011000000000000",--29900
"101010001001101000000001100000000000",--29901
"101111001001110001000011111001001100",--29902
"101111001001100001001100110011001101",--29903
"111110000110001001000001100000000000",--29904
"101111001001110001000011111101100110",--29905
"101111001001100001000110011001100110",--29906
"111110000110010001000010100000000000",--29907
"101110000001111000000001100000000000",--29908
"101110000001111000000010000000000000",--29909
"001001111100000000011111111111011111",--29910
"001011111100000001101111111111011110",--29911
"001001111100000000101111111111011101",--29912
"001001111100000000111111111111011100",--29913
"001001111100000001001111111111011011",--29914
"101000000001111000000000100000000000",--29915
"001001111100000111111111111111011010",--29916
"101001111100010111100000000000100111",--29917
"000111000000000000000110110001101000",--29918
"101001111100000111100000000000100111",--29919
"001101111100000000011111111111011011",--29920
"101010000011101000000001100000000000",--29921
"101111001001110001000011111001001100",--29922
"101111001001100001001100110011001101",--29923
"111110000110001001000001100000000000",--29924
"101111001001110001000011110111001100",--29925
"101111001001100001001100110011001101",--29926
"111110000110000001000010100000000000",--29927
"101000000001111000000000100000000000",--29928
"101110000001111000000001100000000000",--29929
"101110000001111000000010000000000000",--29930
"001101111100000000101111111111011100",--29931
"101001000100000000110000000000000010",--29932
"001111111100000001101111111111011110",--29933
"001101111100000000101111111111011101",--29934
"101001111100010111100000000000100111",--29935
"000111000000000000000110110001101000",--29936
"101001111100000111100000000000100111",--29937
"001101111100000111111111111111011010",--29938
"101001000000000000010000000000000011",--29939
"001101111100000000101111111111011101",--29940
"101001000100000000110000000000000001",--29941
"010111000111000001000000000000000001",--29942
"101001000110010000110000000000000101",--29943
"001111111100000000111111111111011110",--29944
"001101111100000001001111111111011100",--29945
"101000000111111000000001000000000000",--29946
"101000001001111000000001100000000000",--29947
"001001111100000111111111111111011010",--29948
"101001111100010111100000000000100111",--29949
"000111000000000000000110111011001001",--29950
"101001111100000111100000000000100111",--29951
"001101111100000111111111111111011010",--29952
"001101111100000000011111111111011111",--29953
"101001000010010000010000000000000001",--29954
"010111000010000000001111100000000000",--29955
"001101111100000000101111111111011101",--29956
"101001000100000000100000000000000010",--29957
"010111000101000001000000000000000001",--29958
"101001000100010000100000000000000101",--29959
"001101111100000000111111111111011100",--29960
"101001000110000000110000000000000100",--29961
"101010000011101000000001100000000000",--29962
"101111001001110001000011111001001100",--29963
"101111001001100001001100110011001101",--29964
"111110000110001001000001100000000000",--29965
"101111001001110001000011111101100110",--29966
"101111001001100001000110011001100110",--29967
"111110000110010001000001100000000000",--29968
"001001111100000000111111111111011010",--29969
"001001111100000000101111111111011001",--29970
"001001111100000000011111111111011000",--29971
"101001000000000000010000000000000100",--29972
"001001111100000111111111111111010111",--29973
"101001111100010111100000000000101010",--29974
"000111000000000000000110111011001001",--29975
"101001111100000111100000000000101010",--29976
"001101111100000111111111111111010111",--29977
"001101111100000000011111111111011000",--29978
"101001000010010000010000000000000001",--29979
"001101111100000000101111111111011001",--29980
"101001000100000000100000000000000010",--29981
"010111000101000001000000000000000001",--29982
"101001000100010000100000000000000101",--29983
"001101111100000000111111111111011010",--29984
"101001000110000000110000000000000100",--29985
"010111000010000000001111100000000000",--29986
"000101000000000000000111001001010010",--29987
"010111000100000000001111100000000000",--29988
"101110000001111000000001100000000000",--29989
"001001111100000000010000000000000000",--29990
"001001111100000000101111111111111111",--29991
"101001000000000000010000000000000011",--29992
"001001111100000111111111111111111110",--29993
"000111000000000000000111010110110001",--29994
"001101111100000111111111111111111110",--29995
"101000000011111000000001000000000000",--29996
"001101000000000000010000000110101010",--29997
"001001111100000000101111111111111110",--29998
"001001111100000111111111111111111101",--29999
"000111000000000000000111010110101010",--30000
"001101111100000111111111111111111101",--30001
"101000111011111000000001000000000000",--30002
"101001111010000111010000000000000010",--30003
"001001000100000000010000000000000001",--30004
"001101111100000000011111111111111110",--30005
"001001000100000000010000000000000000",--30006
"101000000101111000000000100000000000",--30007
"001101111100000000101111111111111111",--30008
"001101111100000001000000000000000000",--30009
"001000001000000000100000100000000000",--30010
"101001000100010000100000000000000001",--30011
"101000001001111000000000100000000000",--30012
"010111000100000000001111100000000000",--30013
"000101000000000000000111010100100101",--30014
"010111000010000000001111100000000000",--30015
"101001000000000000100000000001111000",--30016
"101110000001111000000001100000000000",--30017
"001001111100000000010000000000000000",--30018
"001001111100000000101111111111111111",--30019
"101001000000000000010000000000000011",--30020
"001001111100000111111111111111111110",--30021
"000111000000000000000111010110110001",--30022
"001101111100000111111111111111111110",--30023
"101000000011111000000001000000000000",--30024
"001101000000000000010000000110101010",--30025
"001001111100000000101111111111111110",--30026
"001001111100000111111111111111111101",--30027
"000111000000000000000111010110101010",--30028
"101000111011111000000001000000000000",--30029
"101001111010000111010000000000000010",--30030
"001001000100000000010000000000000001",--30031
"001101111100000000011111111111111110",--30032
"001001000100000000010000000000000000",--30033
"001101111100000000011111111111111111",--30034
"000111000000000000000111010110101010",--30035
"001101111100000000100000000000000000",--30036
"001001000100000000010000000011111110",--30037
"101001000000000000100000000001110110",--30038
"101001111100010111100000000000000100",--30039
"000111000000000000000111010100100100",--30040
"101001111100000111100000000000000100",--30041
"001101111100000111111111111111111101",--30042
"001101111100000000010000000000000000",--30043
"101001000010010000010000000000000001",--30044
"010111000010000000001111100000000000",--30045
"000101000000000000000111010101000000",--30046
"010111000100000000001111100000000000",--30047
"001100000010000000100001100000000000",--30048
"001001111100000000010000000000000000",--30049
"001001111100000000101111111111111111",--30050
"101000000111111000000000100000000000",--30051
"001001111100000111111111111111111110",--30052
"101001111100010111100000000000000011",--30053
"000111000000000000000000011001101010",--30054
"101001111100000111100000000000000011",--30055
"001101111100000111111111111111111110",--30056
"001101111100000000011111111111111111",--30057
"101001000010010000100000000000000001",--30058
"001101111100000000010000000000000000",--30059
"010111000100000000001111100000000000",--30060
"000101000000000000000111010101100000",--30061
"010111000010000000001111100000000000",--30062
"001101000010000000100000000011111110",--30063
"001001111100000000010000000000000000",--30064
"101000000101111000000000100000000000",--30065
"101001000000000000100000000001110111",--30066
"001001111100000111111111111111111111",--30067
"101001111100010111100000000000000010",--30068
"000111000000000000000111010101011111",--30069
"101001111100000111100000000000000010",--30070
"001101111100000111111111111111111111",--30071
"001101111100000000010000000000000000",--30072
"101001000010010000010000000000000001",--30073
"010111000010000000001111100000000000",--30074
"000101000000000000000111010101101111",--30075
"001001111100000000010000000000000000",--30076
"001001111100000000101111111111111111",--30077
"001011111100000000111111111111111110",--30078
"001011111100000001101111111111111101",--30079
"001011111100000001011111111111111100",--30080
"001011111100000001001111111111111011",--30081
"101001000000000000010000000000000011",--30082
"101110000001111000000001100000000000",--30083
"001001111100000111111111111111111010",--30084
"000111000000000000000111010110110001",--30085
"001101111100000111111111111111111010",--30086
"101000000011111000000001000000000000",--30087
"001101000000000000010000000110101010",--30088
"001001111100000000101111111111111010",--30089
"001001111100000111111111111111111001",--30090
"000111000000000000000111010110101010",--30091
"001101111100000111111111111111111001",--30092
"101000111011111000000001000000000000",--30093
"101001111010000111010000000000000010",--30094
"001001000100000000010000000000000001",--30095
"001101111100000000011111111111111010",--30096
"001001000100000000010000000000000000",--30097
"001111111100000000111111111111111011",--30098
"001011000010000000110000000000000000",--30099
"001111111100000000111111111111111100",--30100
"001011000010000000110000000000000001",--30101
"001111111100000000111111111111111101",--30102
"001011000010000000110000000000000010",--30103
"001001111100000000101111111111111001",--30104
"101000000101111000000000100000000000",--30105
"001001111100000111111111111111111000",--30106
"101001111100010111100000000000001001",--30107
"000111000000000000000000011001101010",--30108
"101001111100000111100000000000001001",--30109
"001101111100000111111111111111111000",--30110
"101000111011111000000000100000000000",--30111
"101001111010000111010000000000000011",--30112
"001111111100000000111111111111111110",--30113
"001011000010000000110000000000000010",--30114
"001101111100000000101111111111111001",--30115
"001001000010000000100000000000000001",--30116
"001101111100000000101111111111111111",--30117
"001001000010000000100000000000000000",--30118
"001101111100000000100000000000000000",--30119
"001001000100000000010000000000000100",--30120
"000100000000000000001111100000000000",--30121
"101000111010000000010001100000000000",--30122
"101000111011111000000000100000000000",--30123
"010100000110000111011111100000000000",--30124
"001001111010000000100000000000000000",--30125
"101001111010000111010000000000000001",--30126
"011100111011000000111111111111111101",--30127
"000100000000000000001111100000000000",--30128
"101000111010000000010001000000000000",--30129
"101000111011111000000000100000000000",--30130
"010100000100000111011111100000000000",--30131
"001011111010000000110000000000000000",--30132
"101001111010000111010000000000000001",--30133
"011100111011000000101111111111111101",--30134
"000100000000000000001111100000000000",--30135
"101111001011110001010100000011001001",--30136
"101111001011100001010000111111011011",--30137
"111110001010011000000010000000000000",--30138
"111110000110001001000010000000000000",--30139
"101110001000110000000010000000000000",--30140
"111110001000001001010010000000000000",--30141
"111110000110010001000001100000000000",--30142
"101111001011110001000100000001001001",--30143
"010110000111000001000000000000000001",--30144
"111110001010010000110001100000000000",--30145
"101111001011110001010011111111001001",--30146
"101111001011110001100011111101001001",--30147
"010110000111000001010000000000011111",--30148
"111110001000010000110001100000000000",--30149
"010110000111000001100000000000010000",--30150
"111110001100010000110001100000000000",--30151
"111110000110001000110010000000000000",--30152
"101111001011110001011011100101001101",--30153
"101111001011100001010110010010110110",--30154
"111110001000001001010010100000000000",--30155
"101111001101110001100011110000001000",--30156
"101111001101100001101000011001100110",--30157
"111110001100000001010010100000000000",--30158
"111110001000001001010010100000000000",--30159
"101111001101110001101011111000101010",--30160
"101111001101100001101010101010101100",--30161
"111110001010000001100010100000000000",--30162
"111110001010001001000010000000000000",--30163
"111110001000000000010010000000000000",--30164
"111110001000001000110001100000000010",--30165
"000100000000000000001111100000000000",--30166
"111110000110001000110001100000000000",--30167
"101111001001110001001011101010110011",--30168
"101111001001100001001000000100000110",--30169
"111110000110001001000010000000000000",--30170
"101111001011110001010011110100101010",--30171
"101111001011100001011010011110001001",--30172
"111110001010000001000010000000000000",--30173
"111110000110001001000010000000000000",--30174
"101111000001110001011011111100000000",--30175
"111110001000000001010010000000000000",--30176
"111110001000001000110001100000000000",--30177
"111110000110000000010001100000000010",--30178
"000100000000000000001111100000000000",--30179
"010110000111000001100000000000010000",--30180
"111110001010010000110001100000000000",--30181
"111110000110001000110010000000000000",--30182
"101111001011110001011011100101001101",--30183
"101111001011100001010110010010110110",--30184
"111110001000001001010010100000000000",--30185
"101111001101110001100011110000001000",--30186
"101111001101100001101000011001100110",--30187
"111110001100000001010010100000000000",--30188
"111110001000001001010010100000000000",--30189
"101111001101110001101011111000101010",--30190
"101111001101100001101010101010101100",--30191
"111110001010000001100010100000000000",--30192
"111110001010001001000010000000000000",--30193
"111110001000000000010010000000000000",--30194
"111110001000001000110001100000000000",--30195
"000100000000000000001111100000000000",--30196
"111110000110001000110001100000000000",--30197
"101111001001110001001011101010110011",--30198
"101111001001100001001000000100000110",--30199
"111110000110001001000010000000000000",--30200
"101111001011110001010011110100101010",--30201
"101111001011100001011010011110001001",--30202
"111110001010000001000010000000000000",--30203
"111110000110001001000010000000000000",--30204
"101111000001110001011011111100000000",--30205
"111110001000000001010010000000000000",--30206
"111110001000001000110001100000000000",--30207
"111110000110000000010001100000000000",--30208
"000100000000000000001111100000000000",--30209
"101111001011110001010100000011001001",--30210
"101111001011100001010000111111011011",--30211
"111110001010011000000010000000000000",--30212
"111110000110001001000010000000000000",--30213
"101110001000110000000010000000000000",--30214
"111110001000001001010010000000000000",--30215
"111110000110010001000001100000000000",--30216
"101111001011110001000100000001001001",--30217
"101111001011110001010011111111001001",--30218
"101111001011110001100011111101001001",--30219
"010110000111000001000000000000100001",--30220
"111110000110010001000001100000000000",--30221
"010110000111000001010000000000000001",--30222
"111110001000010000110001100000000000",--30223
"010110000111000001100000000000001110",--30224
"111110001010010000110001100000000000",--30225
"111110000110001000110001100000000000",--30226
"101111001001110001001011101010110011",--30227
"101111001001100001001000000100000110",--30228
"111110000110001001000010000000000000",--30229
"101111001011110001010011110100101010",--30230
"101111001011100001011010011110001001",--30231
"111110001010000001000010000000000000",--30232
"111110000110001001000010000000000000",--30233
"101111000001110001011011111100000000",--30234
"111110001000000001010010000000000000",--30235
"111110001000001000110001100000000000",--30236
"111110000110000000010001100000000010",--30237
"000100000000000000001111100000000000",--30238
"111110000110001000110010000000000000",--30239
"101111001011110001011011100101001101",--30240
"101111001011100001010110010010110110",--30241
"111110001000001001010010100000000000",--30242
"101111001101110001100011110000001000",--30243
"101111001101100001101000011001100110",--30244
"111110001100000001010010100000000000",--30245
"111110001000001001010010100000000000",--30246
"101111001101110001101011111000101010",--30247
"101111001101100001101010101010101100",--30248
"111110001010000001100010100000000000",--30249
"111110001010001001000010000000000000",--30250
"111110001000000000010010000000000000",--30251
"111110001000001000110001100000000010",--30252
"000100000000000000001111100000000000",--30253
"010110000111000001010000000000000001",--30254
"111110001000010000110001100000000000",--30255
"010110000111000001100000000000001110",--30256
"111110001010010000110001100000000000",--30257
"111110000110001000110001100000000000",--30258
"101111001001110001001011101010110011",--30259
"101111001001100001001000000100000110",--30260
"111110000110001001000010000000000000",--30261
"101111001011110001010011110100101010",--30262
"101111001011100001011010011110001001",--30263
"111110001010000001000010000000000000",--30264
"111110000110001001000010000000000000",--30265
"101111000001110001011011111100000000",--30266
"111110001000000001010010000000000000",--30267
"111110001000001000110001100000000000",--30268
"111110000110000000010001100000000000",--30269
"000100000000000000001111100000000000",--30270
"111110000110001000110010000000000000",--30271
"101111001011110001011011100101001101",--30272
"101111001011100001010110010010110110",--30273
"111110001000001001010010100000000000",--30274
"101111001101110001100011110000001000",--30275
"101111001101100001101000011001100110",--30276
"111110001100000001010010100000000000",--30277
"111110001000001001010010100000000000",--30278
"101111001101110001101011111000101010",--30279
"101111001101100001101010101010101100",--30280
"111110001010000001100010100000000000",--30281
"111110001010001001000010000000000000",--30282
"111110001000000000010010000000000000",--30283
"111110001000001000110001100000000000",--30284
"000100000000000000001111100000000000",--30285
x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000",x"000000000");

begin
  main : process(clk)
  begin
    if rising_edge(clk) then
      if EN = '1' then
        if WE = '1' then
          if din(35 downto 30) /= "100100" then
            mem(conv_integer(addr)) <= din;
          end if;
        else
          inst <= mem(conv_integer(addr));
        end if;
      end if;
    end if;
  end process;
end box;
