-- 固定値の命令メモリ
-- Block RAMを使ったRAM(read-firstだが、実際には書き込みと読み出しは同時には行われない)
-- アドレス幅15bit(形式的に16bitで与える),容量32Kワード
-- fib30にtest1を上書き

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity inst_mem_fixed is
  port (
    clk  : in  std_logic;
    addr : in  std_logic_vector(15 downto 0);
    din  : in  std_logic_vector(31 downto 0);
    inst : out std_logic_vector(31 downto 0);
    EN   : in  std_logic;
    WE   : in  std_logic);
end inst_mem_fixed;

architecture box of inst_mem_fixed is
--  type mem_t is array(0 to 32767) of std_logic_vector(31 downto 0);
  type mem_t is array(0 to 63) of std_logic_vector(31 downto 0);
  signal mem : mem_t := (
    "00011100000000000000100000001111",
"00001100001000000000000000000011",
"00001100001000000000000000000010",
"00001100001000000000000000000001",
"00001100001000000000000000000000",
"11011100000000000000000000001111",
--"10001000000000010000000000011110",
--"00101011110111110000000000000000",
--"10011011110111100000000000000001",
--"01111000000000000000000000001011",
--"10001011110111100000000000000001",
--"00111011110111110000000000000000",
"00001100001000000000000000000011",
"00001100001000000000000000000010",
"00001100001000000000000000000001",
"00001100001000000000000000000000",
"11011100000000000000000000001111",
"10001000000000100000000000000001",
"10011100001000101110000000001101",
"01011011100000000000000000000001",
"01101111111000000000000000001111",
"10011000001000100000000000000001",
"00101011110000010000000000000000",
"10011100010000000000100000001111",
"00101011110111111111111111111111",
"10011011110111100000000000000010",
"01111000000000000000000000001011",
"10001011110111100000000000000010",
"00111011110111111111111111111111",
"00111011110000100000000000000000",
"10011000010000100000000000000010",
"00101011110000011111111111111111",
"10011100010000000000100000001111",
"00101011110111111111111111111110",
"10011011110111100000000000000011",
"01111000000000000000000000001011",
"10001011110111100000000000000011",
"00111011110111111111111111111110",
"00111011110000101111111111111111",
"10011100010000010000100000000000",
"01101111111000000000000000001111",
     x"00000000",--x"00000000",x"00000000",x"00000000",
     x"00000000",x"00000000",x"00000000",x"00000000",
     x"00000000",x"00000000",x"00000000",x"00000000",
     x"00000000",x"00000000",x"00000000",x"00000000",
     x"00000000",x"00000000",x"00000000",x"00000000",
     x"00000000",x"00000000",x"00000000",x"00000000",
     x"00000000",x"00000000",x"00000000",x"00000000",
     x"00000000",x"00000000",x"00000000",x"00000000");


begin
  main : process(clk)
  begin
    if rising_edge(clk) then
      if EN = '1' then
        if WE = '1' then
          mem(conv_integer(addr(5 downto 0))) <= din;
        end if;
        inst <= mem(conv_integer(addr(5 downto 0)));
      end if;
    end if;
  end process;
end box;
